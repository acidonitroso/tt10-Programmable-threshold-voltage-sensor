magic
tech sky130A
magscale 1 2
timestamp 1750413043
<< metal1 >>
rect -2400 13300 -1650 13600
rect -1350 13300 -1344 13600
rect -2400 12900 -2100 13300
rect 4133 11547 4327 11553
rect 3503 11353 4133 11547
rect 4133 11347 4327 11353
rect -2310 10950 2700 11170
rect 3773 10986 5795 11136
rect 3372 10648 4184 10812
rect 4348 10648 4354 10812
rect 3463 9727 4117 9925
rect 4315 9727 4321 9925
rect -1710 9370 2706 9590
rect 5645 9556 5795 10986
rect 3773 9406 5795 9556
rect -1710 8710 -1490 9370
rect 3380 9066 4163 9240
rect 4337 9066 4343 9240
rect -2310 8490 -1490 8710
rect 4117 8359 4315 8365
rect 3471 8161 4117 8359
rect 4117 8155 4315 8161
rect -1700 7800 2716 8020
rect 5645 7976 5795 9406
rect 3773 7967 5797 7976
rect 3773 7826 15199 7967
rect 5645 7817 15199 7826
rect -1700 6210 -1480 7800
rect 3380 7486 4121 7668
rect 4303 7486 4309 7668
rect 3476 6564 4106 6760
rect 4302 6564 4308 6760
rect -2310 5990 -1480 6210
rect -1210 6208 2706 6428
rect 5645 6394 5795 7817
rect 3773 6244 5795 6394
rect -1210 3710 -990 6208
rect 3390 5924 4130 6080
rect 4286 5924 4292 6080
rect 4113 5167 4315 5173
rect 3481 4965 4113 5167
rect 4113 4959 4315 4965
rect -2310 3490 -990 3710
rect -710 4630 2706 4850
rect 5645 4816 5795 6244
rect 3763 4666 5795 4816
rect -710 1210 -490 4630
rect 3374 4322 4118 4502
rect 4298 4322 4304 4502
rect 3481 3419 4123 3609
rect 4313 3419 4319 3609
rect -2310 990 -490 1210
rect -210 3050 2706 3270
rect 5645 3236 5795 4666
rect 3773 3086 5795 3236
rect -210 -1290 10 3050
rect 3378 2754 3772 2910
rect 3928 2754 3934 2910
rect 4125 1997 4283 2003
rect 3473 1839 4125 1997
rect 4125 1833 4283 1839
rect -2310 -1510 10 -1290
rect 290 1470 2706 1690
rect 5645 1656 5795 3086
rect 3773 1506 5795 1656
rect 290 -3790 510 1470
rect 3348 1122 3812 1308
rect 3626 747 3812 1122
rect 3626 555 3812 561
rect 4125 -875 4303 -869
rect 2973 -1053 4125 -875
rect 4125 -1059 4303 -1053
rect -2310 -4010 510 -3790
rect 1090 -1428 2210 -1208
rect 3277 -1243 5477 -1242
rect 5645 -1243 5795 1506
rect 3277 -1392 5795 -1243
rect 5323 -1393 5795 -1392
rect -3150 -6750 -2850 -5150
rect -2400 -6750 -2100 -5800
rect -3156 -7050 -3150 -6750
rect -2850 -7050 -2844 -6750
rect -2400 -7056 -2100 -7050
rect 1090 -7290 1310 -1428
rect 2874 -1760 3360 -1556
rect 3156 -2154 3360 -1760
rect 3156 -2364 3360 -2358
<< via1 >>
rect -1650 13300 -1350 13600
rect 4133 11353 4327 11547
rect 4184 10648 4348 10812
rect 4117 9727 4315 9925
rect 4163 9066 4337 9240
rect 4117 8161 4315 8359
rect 4121 7486 4303 7668
rect 4106 6564 4302 6760
rect 4130 5924 4286 6080
rect 4113 4965 4315 5167
rect 4118 4322 4298 4502
rect 4123 3419 4313 3609
rect 3772 2754 3928 2910
rect 4125 1839 4283 1997
rect 3626 561 3812 747
rect 4125 -1053 4303 -875
rect -3150 -7050 -2850 -6750
rect -2400 -7050 -2100 -6750
rect 3156 -2358 3360 -2154
<< metal2 >>
rect -1650 13600 -1350 13606
rect -1350 13300 -1150 13600
rect -850 13300 -841 13600
rect -1650 13294 -1350 13300
rect 4127 11353 4133 11547
rect 4327 11353 16347 11547
rect 4184 10812 4348 10818
rect 4348 10648 4678 10812
rect 4842 10648 4851 10812
rect 4184 10642 4348 10648
rect 4117 9925 4315 9931
rect 4315 9727 15155 9925
rect 4117 9721 4315 9727
rect 4163 9240 4337 9246
rect 4337 9066 4699 9240
rect 4873 9066 4882 9240
rect 4163 9060 4337 9066
rect 4111 8161 4117 8359
rect 4315 8161 13953 8359
rect 4121 7668 4303 7674
rect 4303 7486 4621 7668
rect 4803 7486 4812 7668
rect 4121 7480 4303 7486
rect 4602 6928 12758 7124
rect 4106 6760 4302 6766
rect 4602 6760 4798 6928
rect 4302 6564 4798 6760
rect 4106 6558 4302 6564
rect 4957 6407 11563 6609
rect 4130 6080 4286 6086
rect 4286 5924 4444 6080
rect 4600 5924 4609 6080
rect 4130 5918 4286 5924
rect 4957 5167 5159 6407
rect 4107 4965 4113 5167
rect 4315 4965 5159 5167
rect 5347 5949 10369 6139
rect 11361 6023 11563 6407
rect 12562 6176 12758 6928
rect 13755 6185 13953 8161
rect 14957 6155 15155 9727
rect 16153 6137 16347 11353
rect 4118 4502 4298 4508
rect 4298 4322 4426 4502
rect 4606 4322 4615 4502
rect 4118 4316 4298 4322
rect 4123 3609 4313 3615
rect 5347 3609 5537 5949
rect 4313 3419 5537 3609
rect 6081 5555 9155 5713
rect 10179 5619 10369 5949
rect 4123 3413 4313 3419
rect 3772 2910 3928 2916
rect 3928 2754 4048 2910
rect 4204 2754 4213 2910
rect 3772 2748 3928 2754
rect 6081 1997 6239 5555
rect 8997 5197 9155 5555
rect 4119 1839 4125 1997
rect 4283 1839 6239 1997
rect 6541 4323 7123 4501
rect 3620 561 3626 747
rect 3812 561 3818 747
rect 3626 200 3812 561
rect 3601 4 3610 200
rect 3806 4 3815 200
rect 6541 1 6719 4323
rect 6541 -158 6721 1
rect 6543 -299 6721 -158
rect 5053 -477 6721 -299
rect 5053 -875 5231 -477
rect 4119 -1053 4125 -875
rect 4303 -1053 5252 -875
rect 3150 -2358 3156 -2154
rect 3360 -2358 3366 -2154
rect 3156 -3034 3360 -2358
rect 3145 -3230 3154 -3034
rect 3350 -3162 3360 -3034
rect 3350 -3230 3359 -3162
rect -3150 -6750 -2850 -6744
rect -2406 -7050 -2400 -6750
rect -2100 -7050 -2094 -6750
rect -3150 -7840 -2850 -7050
rect -2400 -7840 -2100 -7050
<< via2 >>
rect -1150 13300 -850 13600
rect 4678 10648 4842 10812
rect 4699 9066 4873 9240
rect 4621 7486 4803 7668
rect 4444 5924 4600 6080
rect 4426 4322 4606 4502
rect 4048 2754 4204 2910
rect 3610 4 3806 200
rect 3154 -3230 3350 -3034
<< metal3 >>
rect -1155 13600 -845 13605
rect -1155 13300 -1150 13600
rect -850 13300 -50 13600
rect 250 13300 256 13600
rect -1155 13295 -845 13300
rect 4673 10813 4847 10817
rect 4673 10812 7381 10813
rect 4673 10648 4678 10812
rect 4842 10648 7381 10812
rect 4673 10643 7381 10648
rect 4699 10627 7381 10643
rect 4694 9240 6477 9245
rect 4694 9066 4699 9240
rect 4873 9066 6477 9240
rect 4694 9061 6477 9066
rect 4737 9047 6477 9061
rect 4616 7668 4808 7673
rect 4616 7486 4621 7668
rect 4803 7652 4808 7668
rect 4803 7486 5948 7652
rect 4616 7481 5948 7486
rect 4656 7452 5948 7481
rect 4439 6080 5467 6085
rect 4439 5924 4444 6080
rect 4600 5924 5467 6080
rect 4439 5919 5467 5924
rect 4469 5887 5467 5919
rect 4406 4507 4602 4508
rect 4406 4502 4611 4507
rect 4406 4322 4426 4502
rect 4606 4322 4611 4502
rect 4406 4317 4611 4322
rect 4043 2910 4209 2915
rect 4043 2909 4048 2910
rect 4001 2754 4048 2909
rect 4204 2754 4209 2910
rect 4001 2749 4209 2754
rect 3605 200 3811 205
rect 3605 4 3610 200
rect 3806 4 3811 200
rect 3605 -2997 3811 4
rect 4001 -1930 4207 2749
rect 4406 -864 4602 4317
rect 5269 29 5467 5887
rect 5748 1098 5948 7452
rect 6279 2197 6477 9047
rect 7195 4063 7381 10627
rect 4406 -1060 5532 -864
rect 4001 -2136 5517 -1930
rect 3149 -3034 3355 -3029
rect 3149 -3230 3154 -3034
rect 3350 -3230 3355 -3034
rect 3605 -3203 5491 -2997
rect 3149 -4147 3355 -3230
rect 3149 -4353 5507 -4147
<< via3 >>
rect -50 13300 250 13600
<< metal4 >>
rect -51 13600 251 13601
rect -51 13300 -50 13600
rect 250 13300 8686 13600
rect -51 13299 251 13300
rect 1500 11748 1765 13300
rect 1500 11638 2468 11748
rect 1500 10168 1765 11638
rect 1500 10058 2468 10168
rect 1500 8588 1765 10058
rect 1500 8478 2468 8588
rect 1500 7006 1765 8478
rect 1500 6896 2468 7006
rect 1500 5428 1765 6896
rect 1500 5318 2468 5428
rect 1500 3848 1765 5318
rect 1500 3738 2468 3848
rect 1500 2268 1765 3738
rect 1500 2158 2468 2268
rect 1500 -627 1765 2158
rect 1500 -732 1957 -627
rect 1739 -737 1957 -732
rect 3800 -1846 4065 10530
rect 3300 -1956 4065 -1846
rect 3800 -2136 4065 -1956
use partitore_MAGIC  partitore_MAGIC_0
timestamp 1750067613
transform 1 0 -2200 0 1 8350
box -900 -14750 152 5174
use pass_gate_MAGIC  pass_gate_MAGIC_0
timestamp 1749803936
transform 1 0 2518 0 1 1146
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_1
timestamp 1749803936
transform 1 0 2518 0 1 10626
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_2
timestamp 1749803936
transform 1 0 2518 0 1 9046
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_3
timestamp 1749803936
transform 1 0 2518 0 1 7466
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_4
timestamp 1749803936
transform 1 0 2518 0 1 5884
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_5
timestamp 1749803936
transform 1 0 2518 0 1 4306
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_6
timestamp 1749803936
transform 1 0 2518 0 1 2726
box -160 -204 1410 1122
use pass_gate_MAGIC  pass_gate_MAGIC_7
timestamp 1749803936
transform 1 0 2022 0 1 -1752
box -160 -204 1410 1122
<< labels >>
flabel space 3444 11396 3928 11456 0 FreeSans 320 0 960 32 n_d[7]
flabel space 3444 9816 3928 9876 0 FreeSans 320 0 960 32 n_d[6]
flabel space 3444 8236 3928 8296 0 FreeSans 320 0 960 32 n_d[5]
flabel space 3444 6654 3928 6714 0 FreeSans 320 0 960 32 n_d[4]
flabel space 3444 5076 3928 5136 0 FreeSans 320 0 960 32 n_d[3]
flabel space 3444 3496 3928 3556 0 FreeSans 320 0 960 32 n_d[2]
flabel space 3444 1916 3928 1976 0 FreeSans 320 0 960 32 n_d[1]
flabel space 2948 -982 3432 -922 0 FreeSans 320 0 960 32 n_d[0]
flabel space 2849 -1656 3426 -1608 0 FreeSans 320 0 960 32 y_d[0]
flabel space 3345 4402 3922 4450 0 FreeSans 320 0 960 32 y_d[3]
flabel space 3345 5980 3922 6028 0 FreeSans 320 0 960 32 y_d[4]
flabel space 3345 7562 3922 7610 0 FreeSans 320 0 960 32 y_d[5]
flabel space 3345 9142 3922 9190 0 FreeSans 320 0 960 32 y_d[6]
flabel space 3345 10722 3922 10770 0 FreeSans 320 0 960 32 y_d[7]
rlabel metal1 100 10950 2700 11170 1 ete
flabel space 3345 1242 3922 1290 0 FreeSans 320 0 960 32 y_d[1]
flabel space 3345 2822 3922 2870 0 FreeSans 320 0 960 32 y_d[2]
<< end >>
