magic
tech sky130A
magscale 1 2
timestamp 1750694076
<< viali >>
rect -288 2496 -216 2704
rect 308 2502 380 2710
<< metal1 >>
rect -478 5108 580 5560
rect -322 2710 400 2718
rect -322 2704 308 2710
rect -322 2496 -288 2704
rect -216 2502 308 2704
rect 380 2502 400 2710
rect -216 2496 400 2502
rect -322 2480 400 2496
rect -8 1007 202 2480
rect 336 1007 650 1102
rect -991 937 -789 943
rect -8 797 650 1007
rect -991 104 -789 735
rect 336 381 650 797
rect -512 104 -310 106
rect -991 -334 -310 104
rect 336 61 650 67
rect -991 -338 -789 -334
rect -512 -338 -310 -334
<< via1 >>
rect -991 735 -789 937
rect 336 67 650 381
<< metal2 >>
rect -991 1385 -789 1394
rect -991 937 -789 1183
rect -997 735 -991 937
rect -789 735 -783 937
rect 330 67 336 381
rect 650 67 656 381
rect 336 -160 650 -151
<< via2 >>
rect -991 1183 -789 1385
rect 336 67 650 163
rect 336 -151 650 67
<< metal3 >>
rect -991 1883 -789 1889
rect -991 1390 -789 1681
rect -996 1385 -784 1390
rect -996 1183 -991 1385
rect -789 1183 -784 1385
rect -996 1178 -784 1183
rect 331 163 655 168
rect 331 -156 336 163
rect 650 -156 655 163
rect 336 -401 650 -395
<< via3 >>
rect -991 1681 -789 1883
rect 336 -151 650 -81
rect 336 -395 650 -151
<< metal4 >>
rect -991 1884 -789 5705
rect -992 1883 -788 1884
rect -992 1681 -991 1883
rect -789 1681 -788 1883
rect -992 1680 -788 1681
rect 335 -81 651 -80
rect 335 -395 336 -81
rect 650 -395 651 -81
rect 335 -396 651 -395
rect 336 -597 650 -396
use sky130_fd_pr__res_high_po_0p35_MGTKQ5  XR5
timestamp 1749664143
transform 1 0 -403 0 1 2606
box -201 -3102 201 3102
use sky130_fd_pr__res_high_po_0p35_KC2364  XR6
timestamp 1749664143
transform 1 0 497 0 1 3106
box -201 -2612 201 2612
<< end >>
