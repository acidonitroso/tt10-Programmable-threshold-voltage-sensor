magic
tech sky130A
magscale 1 2
timestamp 1750413137
<< viali >>
rect 478 854 630 914
rect 488 -382 640 -322
<< metal1 >>
rect -110 914 684 1004
rect -110 908 478 914
rect -110 722 -14 908
rect 456 854 478 908
rect 630 854 684 914
rect 456 848 684 854
rect 478 846 624 848
rect -110 620 -14 626
rect 66 744 832 816
rect 66 473 138 744
rect 270 706 280 714
rect 354 706 364 714
rect 264 626 274 706
rect 362 626 372 706
rect 526 630 536 714
rect 616 630 626 714
rect 770 630 780 716
rect 876 630 886 716
rect 396 502 406 586
rect 484 502 494 586
rect 650 506 660 584
rect 746 506 756 584
rect 66 408 846 473
rect 66 117 141 408
rect 66 52 652 117
rect 66 51 649 52
rect 66 -212 138 51
rect 520 -56 530 16
rect 598 -56 608 16
rect 424 -178 434 -102
rect 504 -178 514 -102
rect 432 -182 442 -178
rect 496 -182 506 -178
rect 618 -192 628 -112
rect 702 -192 712 -112
rect 66 -276 550 -212
rect 66 -278 138 -276
rect 480 -322 670 -304
rect 1011 -315 1017 -217
rect 1115 -315 1121 -217
rect 480 -355 488 -322
rect 479 -382 488 -355
rect 640 -355 670 -322
rect 1017 -355 1115 -315
rect 640 -382 1115 -355
rect 479 -453 1115 -382
<< via1 >>
rect -110 626 -14 722
rect 280 706 354 714
rect 274 626 362 706
rect 536 630 616 714
rect 780 630 876 716
rect 406 502 484 586
rect 660 506 746 584
rect 530 -56 598 16
rect 434 -178 504 -102
rect 442 -182 496 -178
rect 628 -192 702 -112
rect 1017 -315 1115 -217
<< metal2 >>
rect 280 722 354 724
rect 536 722 616 724
rect 780 722 876 726
rect -116 626 -110 722
rect -14 716 880 722
rect -14 714 780 716
rect -14 706 280 714
rect 354 706 536 714
rect -14 626 274 706
rect 362 630 536 706
rect 616 630 780 714
rect 876 630 880 716
rect 362 626 880 630
rect 274 616 362 626
rect 536 620 616 626
rect 780 620 876 626
rect 406 586 484 596
rect 264 502 406 584
rect 660 584 746 594
rect 484 506 660 584
rect 746 506 1110 584
rect 484 502 1110 506
rect 264 500 1110 502
rect 406 492 484 500
rect 660 496 746 500
rect 1026 30 1110 500
rect 432 16 1110 30
rect 432 -54 530 16
rect 598 -54 1110 16
rect 530 -66 598 -56
rect 434 -102 504 -92
rect 380 -178 434 -104
rect 628 -104 702 -102
rect 504 -112 1115 -104
rect 504 -178 628 -112
rect 380 -182 442 -178
rect 496 -182 628 -178
rect 380 -192 628 -182
rect 702 -192 1115 -112
rect 380 -202 1115 -192
rect 1017 -217 1115 -202
rect 1017 -321 1115 -315
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  sky130_fd_pr__nfet_01v8_lvt_DJ7QE5_0
timestamp 1749574077
transform 1 0 565 0 1 -84
box -263 -310 263 310
use sky130_fd_pr__pfet_01v8_lvt_4QBKD3  sky130_fd_pr__pfet_01v8_lvt_4QBKD3_0
timestamp 1749574077
transform 1 0 573 0 1 615
box -423 -319 423 319
<< end >>
