magic
tech sky130A
magscale 1 2
timestamp 1749663830
<< pwell >>
rect -201 -3592 201 3592
<< psubdiff >>
rect -165 3522 -69 3556
rect 69 3522 165 3556
rect -165 3460 -131 3522
rect 131 3460 165 3522
rect -165 -3522 -131 -3460
rect 131 -3522 165 -3460
rect -165 -3556 -69 -3522
rect 69 -3556 165 -3522
<< psubdiffcont >>
rect -69 3522 69 3556
rect -165 -3460 -131 3460
rect 131 -3460 165 3460
rect -69 -3556 69 -3522
<< xpolycontact >>
rect -35 2994 35 3426
rect -35 -3426 35 -2994
<< ppolyres >>
rect -35 -2994 35 2994
<< locali >>
rect -165 3522 -69 3556
rect 69 3522 165 3556
rect -165 3460 -131 3522
rect 131 3460 165 3522
rect -165 -3522 -131 -3460
rect 131 -3522 165 -3460
rect -165 -3556 -69 -3522
rect 69 -3556 165 -3522
<< viali >>
rect -19 3011 19 3408
rect -19 -3408 19 -3011
<< metal1 >>
rect -25 3408 25 3420
rect -25 3011 -19 3408
rect 19 3011 25 3408
rect -25 2999 25 3011
rect -25 -3011 25 -2999
rect -25 -3408 -19 -3011
rect 19 -3408 25 -3011
rect -25 -3420 25 -3408
<< properties >>
string FIXED_BBOX -148 -3539 148 3539
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 30.1 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 28.616k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
