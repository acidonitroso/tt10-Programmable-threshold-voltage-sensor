magic
tech sky130A
magscale 1 2
timestamp 1750694093
<< metal1 >>
rect 39782 22853 39853 22859
rect 39853 22782 40903 22853
rect 39782 22776 39853 22782
rect 22845 22417 28647 22567
rect 8890 6798 9110 7536
<< via1 >>
rect 39782 22782 39853 22853
<< metal2 >>
rect 27122 23004 27683 23071
rect 39022 22782 39782 22853
rect 39853 22782 39859 22853
rect 19161 20475 19363 20825
rect 20362 20478 20558 20972
rect 21555 20469 21753 20983
rect 22757 20469 22955 20969
rect 23953 20479 24147 20931
rect 16797 19579 16955 19955
rect 17979 19563 18169 20409
rect 14745 18923 15493 19101
rect 4650 7060 4950 7069
rect 5394 6765 5403 7055
rect 5693 6765 5702 7055
rect 4650 6751 4950 6760
<< via2 >>
rect 4650 6760 4950 7060
rect 5403 6765 5693 7055
<< metal3 >>
rect 14995 18447 15181 18849
rect 14079 16471 14277 16995
rect 13548 15414 13748 15898
rect 13069 14641 14007 14839
rect 13132 13540 13990 13736
rect 13109 12464 13985 12670
rect 13085 11397 13977 11603
rect 13067 10247 13985 10453
rect 4645 7060 4955 7065
rect 4645 6760 4650 7060
rect 4950 6760 4955 7060
rect 4645 6755 4955 6760
rect 5398 7055 5698 7060
rect 5398 6765 5403 7055
rect 5693 6765 5698 7055
rect 4650 6518 4950 6755
rect 5398 6517 5698 6765
rect 5393 6219 5399 6517
rect 5697 6219 5703 6517
rect 5398 6218 5698 6219
rect 4650 6212 4950 6218
<< via3 >>
rect 4650 6218 4950 6518
rect 5399 6219 5697 6517
<< metal4 >>
rect 15712 27706 42262 28230
rect 41738 25478 42262 27706
rect 4649 6518 4951 6519
rect 4649 6218 4650 6518
rect 4950 6218 4951 6518
rect 4649 6217 4951 6218
rect 5398 6517 5698 6518
rect 5398 6219 5399 6517
rect 5697 6219 5698 6517
rect 4650 6012 4950 6217
rect 5398 6012 5698 6219
rect 11600 6012 11865 12680
rect 41664 6012 42188 9926
rect 4526 5488 42188 6012
use Matt  Matt_0
timestamp 1750413043
transform 1 0 7800 0 1 14600
box -3156 -7840 16347 13606
use ota  ota_0
timestamp 1750694093
transform 1 0 28462 0 1 19497
box -3790 -9967 13824 6470
<< end >>
