magic
tech sky130A
magscale 1 2
timestamp 1749803936
<< viali >>
rect 471 1040 717 1092
rect 522 -182 708 -122
<< metal1 >>
rect 340 1114 435 1117
rect 340 1112 745 1114
rect 340 1022 355 1112
rect 435 1092 745 1112
rect 435 1040 471 1092
rect 717 1040 745 1092
rect 435 1022 745 1040
rect 510 930 986 990
rect 439 818 449 880
rect 502 818 512 880
rect 690 816 700 878
rect 760 816 770 878
rect 926 830 986 930
rect 926 770 1410 830
rect 559 706 569 767
rect 633 706 643 767
rect 926 670 986 770
rect 510 610 986 670
rect 141 539 151 551
rect -56 326 151 539
rect 141 324 151 326
rect 238 324 248 551
rect 1000 340 1010 530
rect 1100 510 1110 530
rect 1100 360 1405 510
rect 1100 340 1110 360
rect 565 243 876 291
rect 511 69 521 159
rect 579 69 589 159
rect 626 69 636 159
rect 689 69 699 159
rect 827 144 875 243
rect 827 96 1224 144
rect 827 -27 875 96
rect 564 -75 875 -27
rect 483 -122 793 -104
rect 483 -182 522 -122
rect 708 -182 793 -122
rect 483 -194 793 -182
rect 873 -194 888 -104
rect 483 -196 888 -194
rect 793 -199 888 -196
<< via1 >>
rect 355 1022 435 1112
rect 449 818 502 880
rect 700 816 760 878
rect 569 706 633 767
rect 151 324 238 551
rect 1010 340 1100 530
rect 521 69 579 159
rect 636 69 689 159
rect 793 -194 873 -104
<< metal2 >>
rect 225 1112 435 1122
rect 225 1022 245 1112
rect 325 1022 355 1112
rect 225 1012 435 1022
rect 449 889 502 890
rect 420 885 1110 889
rect 420 880 1115 885
rect 420 818 449 880
rect 502 878 1115 880
rect 502 818 700 878
rect 420 816 700 818
rect 760 816 1115 878
rect 420 808 1115 816
rect 700 806 760 808
rect 132 767 650 780
rect 132 706 569 767
rect 633 706 650 767
rect 132 700 650 706
rect 132 551 258 700
rect 569 696 633 700
rect 132 324 151 551
rect 238 324 258 551
rect 132 177 258 324
rect 985 530 1115 808
rect 985 340 1010 530
rect 1100 340 1115 530
rect 985 179 1115 340
rect 132 159 589 177
rect 132 69 521 159
rect 579 69 589 159
rect 132 51 589 69
rect 628 159 1115 179
rect 628 69 636 159
rect 689 69 1115 159
rect 628 49 1115 69
rect 793 -104 1003 -94
rect 873 -194 903 -104
rect 983 -194 1003 -104
rect 793 -204 1003 -194
<< via2 >>
rect 245 1022 325 1112
rect 903 -194 983 -104
<< metal3 >>
rect 125 1117 295 1122
rect 125 1112 335 1117
rect 125 1022 135 1112
rect 215 1022 245 1112
rect 325 1022 335 1112
rect 125 1017 335 1022
rect 125 1012 295 1017
rect 933 -99 1103 -94
rect 893 -104 1103 -99
rect 893 -194 903 -104
rect 983 -194 1013 -104
rect 1093 -194 1103 -104
rect 893 -199 1103 -194
rect 933 -204 1103 -199
<< via3 >>
rect 135 1022 215 1112
rect 1013 -194 1093 -104
<< metal4 >>
rect -160 1113 195 1122
rect -160 1112 216 1113
rect -160 1022 135 1112
rect 215 1022 216 1112
rect -160 1021 216 1022
rect -160 1012 195 1021
rect 1033 -103 1388 -94
rect 1012 -104 1388 -103
rect 1012 -194 1013 -104
rect 1093 -194 1388 -104
rect 1012 -195 1388 -194
rect 1033 -204 1388 -195
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM11
timestamp 1749574077
transform -1 0 611 0 -1 110
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM23
timestamp 1749567790
transform -1 0 605 0 -1 799
box -295 -319 295 319
<< end >>
