magic
tech sky130A
magscale 1 2
timestamp 1750694093
<< viali >>
rect -172 3590 -94 3800
rect 386 3596 464 3806
<< metal1 >>
rect -364 6080 660 6546
rect -206 3806 492 3814
rect -206 3800 386 3806
rect -206 3590 -172 3800
rect -94 3596 386 3800
rect 464 3596 492 3806
rect -94 3590 492 3596
rect -206 3572 492 3590
rect -798 1816 -566 1822
rect -798 1094 -566 1584
rect -806 596 -172 1094
rect 98 902 302 3572
rect 406 902 752 1092
rect 98 698 752 902
rect -798 594 -566 596
rect -406 594 -174 596
rect 406 407 752 698
rect 406 55 752 61
<< via1 >>
rect -798 1584 -566 1816
rect 406 61 752 407
<< metal2 >>
rect -798 2286 -566 2295
rect -798 1816 -566 2054
rect -804 1584 -798 1816
rect -566 1584 -560 1816
rect 400 61 406 407
rect 752 61 758 407
rect 406 -198 752 -189
<< via2 >>
rect -798 2054 -566 2286
rect 406 61 752 157
rect 406 -189 752 61
<< metal3 >>
rect -798 2864 -566 2870
rect -798 2291 -566 2632
rect -803 2286 -561 2291
rect -803 2054 -798 2286
rect -566 2054 -561 2286
rect -803 2049 -561 2054
rect 401 157 757 162
rect 401 -194 406 157
rect 752 -194 757 157
rect 406 -409 752 -403
<< via3 >>
rect -798 2632 -566 2864
rect 406 -189 752 -57
rect 406 -403 752 -189
<< metal4 >>
rect -798 2865 -566 6668
rect -799 2864 -565 2865
rect -799 2632 -798 2864
rect -566 2632 -565 2864
rect -799 2631 -565 2632
rect 405 -57 753 -56
rect 405 -403 406 -57
rect 752 -403 753 -57
rect 405 -404 753 -403
rect 406 -601 752 -404
use sky130_fd_pr__res_high_po_0p35_MGTKQ5  XR2
timestamp 1749664143
transform 1 0 -285 0 1 3598
box -201 -3102 201 3102
use sky130_fd_pr__res_high_po_0p35_MGTKQ5  XR3
timestamp 1749664143
transform 1 0 579 0 1 3596
box -201 -3102 201 3102
<< end >>
