magic
tech sky130A
magscale 1 2
timestamp 1750669323
<< metal1 >>
rect 2180 41852 26560 41908
rect 26616 41852 26622 41908
rect 2180 20856 2236 41852
rect 2922 41076 2978 41078
rect 2922 41020 27102 41076
rect 27158 41020 27190 41076
rect 2922 24168 2978 41020
rect 5780 40014 27788 40022
rect 5780 39966 27656 40014
rect 5780 39614 5836 39966
rect 27650 39958 27656 39966
rect 27712 39966 27788 40014
rect 27712 39958 27718 39966
rect 5774 39558 5780 39614
rect 5836 39558 5842 39614
rect 2922 24106 2978 24112
rect 2180 20794 2236 20800
rect 4036 950 4256 35178
rect 20034 1494 20105 3244
rect 20034 1423 26571 1494
rect 4036 730 19134 950
rect 19354 730 19360 950
rect 26500 899 26571 1423
rect 26496 839 26571 899
rect 26496 802 26567 839
rect 26496 725 26567 731
<< via1 >>
rect 26560 41852 26616 41908
rect 27102 41020 27158 41076
rect 27656 39958 27712 40014
rect 5780 39558 5836 39614
rect 2922 24112 2978 24168
rect 2180 20800 2236 20856
rect 19134 730 19354 950
rect 26496 731 26567 802
<< metal2 >>
rect 26558 44696 26618 44705
rect 27654 44704 27714 44713
rect 26558 44627 26618 44636
rect 27100 44692 27160 44701
rect 27654 44635 27714 44644
rect 26560 41908 26616 44627
rect 27100 44623 27160 44632
rect 26560 41798 26616 41852
rect 27102 41076 27158 44623
rect 27102 41014 27158 41020
rect 27656 40014 27712 44635
rect 27656 39952 27712 39958
rect 5780 39614 5836 39620
rect 5780 27424 5836 39558
rect 16161 28465 16339 28753
rect 15379 28287 16339 28465
rect 15369 27113 16975 27271
rect 15371 25899 16991 26089
rect 15367 24705 17915 24907
rect 2916 24112 2922 24168
rect 2978 24112 5826 24168
rect 15370 23510 17912 23706
rect 15585 22315 17919 22513
rect 15563 21113 17905 21311
rect 2174 20800 2180 20856
rect 2236 20800 5826 20856
rect 15557 19921 17911 20115
rect 20242 16879 26509 16946
rect 26442 2494 26509 16879
rect 26442 2427 30495 2494
rect 30428 1676 30495 2427
rect 30428 1600 30495 1609
rect 19134 950 19354 956
rect 19354 730 20088 950
rect 20308 730 20317 950
rect 26490 731 26496 802
rect 26567 731 26573 802
rect 19134 724 19354 730
rect 26496 638 26567 731
rect 26496 558 26567 567
<< via2 >>
rect 26558 44636 26618 44696
rect 27100 44632 27160 44692
rect 27654 44644 27714 44704
rect 30428 1609 30495 1676
rect 20088 730 20308 950
rect 26496 567 26567 638
<< metal3 >>
rect 27098 44866 27162 44872
rect 26556 44858 26620 44864
rect 27098 44796 27162 44802
rect 27652 44866 27716 44872
rect 27652 44796 27716 44802
rect 26556 44788 26620 44794
rect 26558 44701 26618 44788
rect 26553 44696 26623 44701
rect 27100 44697 27160 44796
rect 27654 44709 27714 44796
rect 27649 44704 27719 44709
rect 26553 44636 26558 44696
rect 26618 44636 26623 44696
rect 26553 44631 26623 44636
rect 27095 44692 27165 44697
rect 27095 44632 27100 44692
rect 27160 44632 27165 44692
rect 27649 44644 27654 44704
rect 27714 44644 27719 44704
rect 27649 44639 27719 44644
rect 27095 44627 27165 44632
rect 1537 41764 1935 41769
rect 186 41364 192 41764
rect 592 41763 1936 41764
rect 592 41365 1537 41763
rect 1935 41365 1936 41763
rect 592 41364 1936 41365
rect 1537 41359 1935 41364
rect 7485 29981 7691 30289
rect 6823 29775 7691 29981
rect 6823 28921 7029 29775
rect 8635 29711 8841 30297
rect 7909 29505 8841 29711
rect 7909 28929 8115 29505
rect 9702 29467 9908 30289
rect 8999 29261 9908 29467
rect 8999 28899 9205 29261
rect 10778 29108 10974 30274
rect 10024 28912 10974 29108
rect 11879 29101 12077 30259
rect 12652 29106 12852 30520
rect 13709 29113 13907 29989
rect 11211 28903 12077 29101
rect 12308 28906 12852 29106
rect 13391 28915 13907 29113
rect 14477 28887 15871 29073
rect 30423 1676 30500 1681
rect 30423 1609 30428 1676
rect 30495 1609 30500 1676
rect 30423 1604 30500 1609
rect 30428 1174 30495 1604
rect 30428 1101 30495 1107
rect 20083 950 20313 955
rect 20083 730 20088 950
rect 20308 730 21616 950
rect 21836 730 21842 950
rect 20083 725 20313 730
rect 26491 638 26572 643
rect 26491 567 26496 638
rect 26567 567 26572 638
rect 26491 562 26572 567
rect 26496 470 26567 562
rect 26496 393 26567 399
<< via3 >>
rect 26556 44794 26620 44858
rect 27098 44802 27162 44866
rect 27652 44802 27716 44866
rect 192 41364 592 41764
rect 1537 41365 1935 41763
rect 30428 1107 30495 1174
rect 21616 730 21836 950
rect 26496 399 26567 470
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 44152 18338 45152
rect 18830 44152 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44859 26618 45152
rect 27110 45074 27170 45152
rect 27662 45078 27722 45152
rect 27100 44952 27170 45074
rect 27654 44952 27722 45078
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27100 44867 27160 44952
rect 27654 44867 27714 44952
rect 27097 44866 27163 44867
rect 26555 44858 26621 44859
rect 26555 44794 26556 44858
rect 26620 44794 26621 44858
rect 27097 44802 27098 44866
rect 27162 44802 27163 44866
rect 27097 44801 27163 44802
rect 27651 44866 27717 44867
rect 27651 44802 27652 44866
rect 27716 44802 27717 44866
rect 27651 44801 27717 44802
rect 26555 44793 26621 44794
rect 200 41765 600 44152
rect 191 41764 600 41765
rect 191 41364 192 41764
rect 592 41364 600 41764
rect 191 41363 600 41364
rect 200 1000 600 41363
rect 800 43752 19276 44152
rect 800 37180 1200 43752
rect 1536 41763 26978 41764
rect 1536 41365 1537 41763
rect 1935 41365 26978 41763
rect 1536 41364 26978 41365
rect 800 36656 3250 37180
rect 800 1000 1200 36656
rect 26578 27180 26978 41364
rect 25166 26780 26978 27180
rect 2848 24850 7728 25170
rect 13534 24862 25254 25182
rect 30427 1174 30496 1175
rect 30427 1107 30428 1174
rect 30495 1107 30496 1174
rect 30427 1106 30496 1107
rect 21615 950 21837 951
rect 21615 730 21616 950
rect 21836 730 22812 950
rect 21615 729 21837 730
rect 22592 200 22812 730
rect 26495 470 26568 471
rect 26495 399 26496 470
rect 26567 399 26568 470
rect 26495 398 26568 399
rect 26496 200 26567 398
rect 30428 200 30495 1106
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22592 0 22814 200
rect 26496 123 26678 200
rect 26498 0 26678 123
rect 30362 0 30542 200
rect 22592 -6 22812 0
use analog  analog_0
timestamp 1750431682
transform 0 1 -2748 -1 0 44076
box 4526 5488 42286 28230
use decoder_p  decoder_p_0
timestamp 1750432038
transform 0 1 5770 -1 0 29154
box 0 0 9186 10000
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
