magic
tech sky130A
magscale 1 2
timestamp 1749567790
<< error_p >>
rect -95 181 -33 187
rect 33 181 95 187
rect -95 147 -83 181
rect 33 147 45 181
rect -95 141 -33 147
rect 33 141 95 147
rect -95 -147 -33 -141
rect 33 -147 95 -141
rect -95 -181 -83 -147
rect 33 -181 45 -147
rect -95 -187 -33 -181
rect 33 -187 95 -181
<< nwell >>
rect -295 -319 295 319
<< pmoslvt >>
rect -99 -100 -29 100
rect 29 -100 99 100
<< pdiff >>
rect -157 88 -99 100
rect -157 -88 -145 88
rect -111 -88 -99 88
rect -157 -100 -99 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 99 88 157 100
rect 99 -88 111 88
rect 145 -88 157 88
rect 99 -100 157 -88
<< pdiffc >>
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
<< nsubdiff >>
rect -259 249 -163 283
rect 163 249 259 283
rect -259 187 -225 249
rect 225 187 259 249
rect -259 -249 -225 -187
rect 225 -249 259 -187
rect -259 -283 -163 -249
rect 163 -283 259 -249
<< nsubdiffcont >>
rect -163 249 163 283
rect -259 -187 -225 187
rect 225 -187 259 187
rect -163 -283 163 -249
<< poly >>
rect -99 181 -29 197
rect -99 147 -83 181
rect -45 147 -29 181
rect -99 100 -29 147
rect 29 181 99 197
rect 29 147 45 181
rect 83 147 99 181
rect 29 100 99 147
rect -99 -147 -29 -100
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect -99 -197 -29 -181
rect 29 -147 99 -100
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 29 -197 99 -181
<< polycont >>
rect -83 147 -45 181
rect 45 147 83 181
rect -83 -181 -45 -147
rect 45 -181 83 -147
<< locali >>
rect -259 249 -163 283
rect 163 249 259 283
rect -259 187 -225 249
rect 225 187 259 249
rect -99 147 -83 181
rect -45 147 -29 181
rect 29 147 45 181
rect 83 147 99 181
rect -145 88 -111 104
rect -145 -104 -111 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 111 88 145 104
rect 111 -104 145 -88
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 83 -181 99 -147
rect -259 -249 -225 -187
rect 225 -249 259 -187
rect -259 -283 -163 -249
rect 163 -283 259 -249
<< viali >>
rect -83 147 -45 181
rect 45 147 83 181
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect -83 -181 -45 -147
rect 45 -181 83 -147
<< metal1 >>
rect -95 181 -33 187
rect -95 147 -83 181
rect -45 147 -33 181
rect -95 141 -33 147
rect 33 181 95 187
rect 33 147 45 181
rect 83 147 95 181
rect 33 141 95 147
rect -151 88 -105 100
rect -151 -88 -145 88
rect -111 -88 -105 88
rect -151 -100 -105 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 105 88 151 100
rect 105 -88 111 88
rect 145 -88 151 88
rect 105 -100 151 -88
rect -95 -147 -33 -141
rect -95 -181 -83 -147
rect -45 -181 -33 -147
rect -95 -187 -33 -181
rect 33 -147 95 -141
rect 33 -181 45 -147
rect 83 -181 95 -147
rect 33 -187 95 -181
<< properties >>
string FIXED_BBOX -242 -266 242 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
