magic
tech sky130A
magscale 1 2
timestamp 1750694093
<< metal1 >>
rect 4427 5263 4502 5269
rect 4427 4946 4502 5188
rect 6178 5254 6255 5260
rect 6178 4942 6255 5177
rect 9906 5166 10018 5172
rect 7202 5155 7277 5161
rect 7202 4071 7277 5080
rect 8522 5150 8634 5156
rect 8522 4006 8634 5038
rect 9906 4038 10018 5054
rect 6570 3438 6641 3444
rect 6641 3367 6975 3438
rect 7785 3375 7851 3381
rect 6570 3361 6641 3367
rect 7851 3309 8103 3375
rect 9164 3344 9235 3350
rect 7785 3303 7851 3309
rect 9235 3273 9501 3344
rect 9164 3267 9235 3273
rect -854 2994 478 3054
rect 4426 1466 4509 1745
rect 6194 1546 6277 1745
rect 7258 1698 7341 2515
rect 7258 1609 7341 1615
rect 8526 1716 8638 2634
rect 8526 1598 8638 1604
rect 9922 1710 10034 2718
rect 9922 1592 10034 1598
rect 4420 1383 4426 1466
rect 4509 1383 4515 1466
rect 5018 1412 5024 1489
rect 5101 1412 5107 1489
rect 6194 1457 6277 1463
rect 5024 37 5101 1412
rect 5136 1292 5142 1364
rect 5214 1292 5220 1364
rect 5429 1303 5435 1377
rect 5509 1303 5515 1377
rect 4484 -40 5101 37
rect 5142 56 5214 1292
rect 5435 987 5509 1303
rect 5435 913 10013 987
rect 5142 -16 7300 56
rect 1937 -469 1999 -463
rect -788 -1452 -782 -1392
rect -722 -1452 -716 -1392
rect -782 -2008 -722 -1452
rect 1937 -2013 1999 -531
rect 4484 -1930 4561 -40
rect 7228 -2004 7300 -16
rect 9939 -2009 10013 913
<< via1 >>
rect 4427 5188 4502 5263
rect 6178 5177 6255 5254
rect 7202 5080 7277 5155
rect 8522 5038 8634 5150
rect 9906 5054 10018 5166
rect 6570 3367 6641 3438
rect 7785 3309 7851 3375
rect 9164 3273 9235 3344
rect 7258 1615 7341 1698
rect 8526 1604 8638 1716
rect 9922 1598 10034 1710
rect 4426 1383 4509 1466
rect 5024 1412 5101 1489
rect 6194 1463 6277 1546
rect 5142 1292 5214 1364
rect 5435 1303 5509 1377
rect 1937 -531 1999 -469
rect -782 -1452 -722 -1392
<< metal2 >>
rect 4427 5425 4502 5434
rect 4427 5263 4502 5350
rect 6178 5416 6255 5425
rect 9906 5374 10018 5383
rect 8522 5362 8634 5371
rect 4421 5188 4427 5263
rect 4502 5188 4508 5263
rect 6178 5254 6255 5339
rect 7202 5341 7277 5350
rect 6172 5177 6178 5254
rect 6255 5177 6261 5254
rect 7202 5155 7277 5266
rect 7196 5080 7202 5155
rect 7277 5080 7283 5155
rect 8522 5150 8634 5250
rect 9906 5166 10018 5262
rect 8516 5038 8522 5150
rect 8634 5038 8640 5150
rect 9900 5054 9906 5166
rect 10018 5054 10024 5166
rect -151 4738 -142 4798
rect -82 4738 468 4798
rect 3596 4458 3659 4462
rect 3591 4453 4462 4458
rect 3591 4390 3596 4453
rect 3659 4390 4462 4453
rect 3591 4385 4462 4390
rect 3596 4381 3659 4385
rect 6338 3934 6401 3938
rect 3438 3861 3573 3934
rect 3646 3861 3655 3934
rect 6218 3929 6406 3934
rect 6218 3866 6338 3929
rect 6401 3866 6406 3929
rect 6218 3861 6406 3866
rect 6338 3857 6401 3861
rect -877 3506 519 3573
rect 6196 3367 6570 3438
rect 6641 3367 6647 3438
rect 7637 3309 7785 3375
rect 7851 3309 7857 3375
rect 9016 3273 9164 3344
rect 9235 3273 9241 3344
rect 10412 3278 11113 3349
rect 3458 3004 3701 3086
rect 3783 3004 3792 3086
rect 3670 2607 4484 2612
rect 3666 2533 3675 2607
rect 3749 2533 4484 2607
rect 3670 2528 4484 2533
rect 6213 2566 6419 2571
rect 6213 2494 6342 2566
rect 6414 2494 6423 2566
rect 6213 2489 6419 2494
rect 378 -469 440 1975
rect 7252 1615 7258 1698
rect 7341 1615 7347 1698
rect 5024 1489 5101 1590
rect 7258 1550 7341 1615
rect 8520 1604 8526 1716
rect 8638 1604 8644 1716
rect 4426 1466 4509 1472
rect 6188 1463 6194 1546
rect 6277 1463 6283 1546
rect 5435 1448 5509 1453
rect 5142 1439 5214 1444
rect 5024 1406 5101 1412
rect 4426 1284 4509 1383
rect 5138 1377 5147 1439
rect 5209 1377 5218 1439
rect 5431 1384 5440 1448
rect 5504 1384 5513 1448
rect 5435 1377 5509 1384
rect 5142 1364 5214 1377
rect 5435 1297 5509 1303
rect 6194 1350 6277 1463
rect 7258 1458 7341 1467
rect 8526 1568 8638 1604
rect 9916 1598 9922 1710
rect 10034 1598 10040 1710
rect 8526 1447 8638 1456
rect 9922 1568 10034 1598
rect 9922 1447 10034 1456
rect 5142 1286 5214 1292
rect 6194 1258 6277 1267
rect 4426 1192 4509 1201
rect -780 -478 -724 -471
rect -782 -480 -722 -478
rect -782 -536 -780 -480
rect -724 -536 -722 -480
rect 378 -531 1937 -469
rect 1999 -531 2005 -469
rect -782 -1392 -722 -536
rect -782 -1458 -722 -1452
<< via2 >>
rect 4427 5350 4502 5425
rect 6178 5339 6255 5416
rect 7202 5266 7277 5341
rect 8522 5250 8634 5362
rect 9906 5262 10018 5374
rect -142 4738 -82 4798
rect 3596 4390 3659 4453
rect 3573 3861 3646 3934
rect 6338 3866 6401 3929
rect 3701 3004 3783 3086
rect 3675 2533 3749 2607
rect 6342 2494 6414 2566
rect 7258 1467 7341 1550
rect 5147 1377 5209 1439
rect 5440 1384 5504 1448
rect 8526 1456 8638 1568
rect 9922 1456 10034 1568
rect 4426 1201 4509 1284
rect 6194 1267 6277 1350
rect -780 -536 -724 -480
<< metal3 >>
rect 6178 5594 6255 5600
rect 4427 5563 4502 5569
rect 4427 5430 4502 5488
rect 9906 5536 10018 5542
rect 4422 5425 4507 5430
rect 4422 5350 4427 5425
rect 4502 5350 4507 5425
rect 6178 5421 6255 5517
rect 8522 5528 8634 5534
rect 7202 5493 7277 5499
rect 4422 5345 4507 5350
rect 6173 5416 6260 5421
rect 6173 5339 6178 5416
rect 6255 5339 6260 5416
rect 7202 5346 7277 5418
rect 8522 5367 8634 5416
rect 9906 5379 10018 5424
rect 9901 5374 10023 5379
rect 8517 5362 8639 5367
rect 6173 5334 6260 5339
rect 7197 5341 7282 5346
rect 7197 5266 7202 5341
rect 7277 5266 7282 5341
rect 7197 5261 7282 5266
rect 8517 5250 8522 5362
rect 8634 5250 8639 5362
rect 9901 5262 9906 5374
rect 10018 5262 10023 5374
rect 9901 5257 10023 5262
rect 8517 5245 8639 5250
rect -147 4798 -77 4803
rect -147 4738 -142 4798
rect -82 4738 -77 4798
rect -147 4733 -77 4738
rect -785 -478 -719 -475
rect -142 -478 -82 4733
rect 3426 4453 3664 4458
rect 3426 4390 3596 4453
rect 3659 4390 3664 4453
rect 3426 4385 3664 4390
rect 3568 3934 3651 3939
rect 3568 3861 3573 3934
rect 3646 3929 6406 3934
rect 3646 3866 6338 3929
rect 6401 3866 6406 3929
rect 3646 3861 6406 3866
rect 3568 3856 3651 3861
rect 3696 3086 3788 3091
rect 3696 3004 3701 3086
rect 3783 3004 6419 3086
rect 3696 2999 3788 3004
rect 3457 2607 3754 2612
rect 3457 2533 3675 2607
rect 3749 2533 3754 2607
rect 3457 2528 3754 2533
rect 6337 2566 6419 3004
rect 6337 2494 6342 2566
rect 6414 2494 6419 2566
rect 6337 2489 6419 2494
rect 8521 1568 8643 1573
rect 7253 1550 7346 1555
rect 5142 1439 5214 1538
rect 5142 1377 5147 1439
rect 5209 1377 5214 1439
rect 5435 1448 5509 1533
rect 7253 1467 7258 1550
rect 7341 1467 7346 1550
rect 7253 1462 7346 1467
rect 5435 1384 5440 1448
rect 5504 1384 5509 1448
rect 5435 1379 5509 1384
rect 7258 1418 7341 1462
rect 8521 1456 8526 1568
rect 8638 1456 8643 1568
rect 8521 1451 8643 1456
rect 9917 1568 10039 1573
rect 9917 1456 9922 1568
rect 10034 1456 10039 1568
rect 9917 1451 10039 1456
rect 5142 1372 5214 1377
rect 6189 1350 6282 1355
rect 4421 1284 4514 1289
rect 4421 1201 4426 1284
rect 4509 1201 4514 1284
rect 6189 1267 6194 1350
rect 6277 1267 6282 1350
rect 7258 1329 7341 1335
rect 8526 1426 8638 1451
rect 8526 1308 8638 1314
rect 9922 1428 10034 1451
rect 9922 1310 10034 1316
rect 6189 1262 6282 1267
rect 4421 1196 4514 1201
rect 4426 1112 4509 1196
rect 6194 1192 6277 1262
rect 4420 1029 4426 1112
rect 4509 1029 4515 1112
rect 6194 1103 6277 1109
rect -785 -480 -82 -478
rect -785 -536 -780 -480
rect -724 -536 -82 -480
rect -785 -538 -82 -536
rect -785 -541 -719 -538
<< via3 >>
rect 4427 5488 4502 5563
rect 6178 5517 6255 5594
rect 7202 5418 7277 5493
rect 8522 5416 8634 5528
rect 9906 5424 10018 5536
rect 7258 1335 7341 1418
rect 8526 1314 8638 1426
rect 9922 1316 10034 1428
rect 4426 1029 4509 1112
rect 6194 1109 6277 1192
<< metal4 >>
rect 9906 6372 10018 6380
rect -86 5848 13824 6372
rect 4427 5564 4502 5848
rect 6178 5595 6255 5848
rect 6177 5594 6256 5595
rect 4426 5563 4503 5564
rect 4426 5488 4427 5563
rect 4502 5488 4503 5563
rect 6177 5517 6178 5594
rect 6255 5517 6256 5594
rect 6177 5516 6256 5517
rect 7202 5494 7277 5848
rect 8522 5529 8634 5848
rect 9906 5537 10018 5848
rect 9905 5536 10019 5537
rect 8521 5528 8635 5529
rect 4426 5487 4503 5488
rect 7201 5493 7278 5494
rect 7201 5418 7202 5493
rect 7277 5418 7278 5493
rect 7201 5417 7278 5418
rect 8521 5416 8522 5528
rect 8634 5416 8635 5528
rect 9905 5424 9906 5536
rect 10018 5424 10019 5536
rect 9905 5423 10019 5424
rect 8521 5415 8635 5416
rect 9921 1428 10035 1429
rect 8525 1426 8639 1427
rect 7257 1418 7342 1419
rect 7257 1335 7258 1418
rect 7341 1335 7342 1418
rect 7257 1334 7342 1335
rect 6193 1192 6278 1193
rect 4425 1112 4510 1113
rect 4425 1029 4426 1112
rect 4509 1029 4510 1112
rect 6193 1109 6194 1192
rect 6277 1109 6278 1192
rect 6193 1108 6278 1109
rect 4425 1028 4510 1029
rect -3790 848 -3266 862
rect 4426 848 4509 1028
rect 6194 848 6277 1108
rect 7258 848 7341 1334
rect 8525 1314 8526 1426
rect 8638 1314 8639 1426
rect 9921 1316 9922 1428
rect 10034 1316 10035 1428
rect 9921 1315 10035 1316
rect 8525 1313 8639 1314
rect 8526 848 8638 1313
rect 9922 848 10034 1315
rect -3790 324 10288 848
rect -3790 -9378 -3266 324
rect 13300 -740 13824 5848
rect -2093 -1258 13824 -740
rect -2093 -1264 13504 -1258
rect -1771 -2091 -1549 -1264
rect 918 -2079 1117 -1264
rect 3586 -1882 3806 -1264
rect 6193 -2373 6395 -1264
rect 9122 -2208 9354 -1264
rect -538 -9378 -228 -6700
rect 2172 -9378 2502 -7942
rect 7532 -9378 7826 -7970
rect 10330 -9378 10676 -8988
rect -3790 -9902 13766 -9378
use carico  carico_0
timestamp 1750693988
transform 1 0 3528 0 1 5012
box 890 -3500 2755 17
use ingresso_ota  ingresso_ota_0
timestamp 1750693945
transform 1 0 -289 0 1 4906
box 501 -4682 3830 1564
use inverter_fine  inverter_fine_0
timestamp 1750413137
transform 1 0 8016 0 1 3076
box -116 -453 1121 1004
use inverter_fine  inverter_fine_1
timestamp 1750413137
transform 1 0 9412 0 1 3082
box -116 -453 1121 1004
use inverter_primo  inverter_primo_0
timestamp 1750416658
transform 1 0 6690 0 1 1784
box 138 698 1016 2318
use vb1_part  vb1_part_0
timestamp 1750694058
transform 1 0 4684 0 1 -9367
box -1104 -600 502 7902
use vb2_part  vb2_part_0
timestamp 1750694076
transform 1 0 7184 0 1 -7427
box -997 -597 698 5718
use vb3_part  vb3_part_0
timestamp 1750694093
transform 1 0 9920 0 1 -8432
box -806 -601 780 6700
use vmirnmos  vmirnmos_0
timestamp 1750694016
transform 1 0 -1324 0 1 -9446
box -458 530 1154 7731
use vmirpmos  vmirpmos_0
timestamp 1750694029
transform 1 0 1312 0 1 -8481
box -400 499 1218 6751
<< end >>
