magic
tech sky130A
magscale 1 2
timestamp 1750063742
<< pwell >>
rect -201 -1212 201 1212
<< psubdiff >>
rect -165 1142 -69 1176
rect 69 1142 165 1176
rect -165 1080 -131 1142
rect 131 1080 165 1142
rect -165 -1142 -131 -1080
rect 131 -1142 165 -1080
rect -165 -1176 -69 -1142
rect 69 -1176 165 -1142
<< psubdiffcont >>
rect -69 1142 69 1176
rect -165 -1080 -131 1080
rect 131 -1080 165 1080
rect -69 -1176 69 -1142
<< xpolycontact >>
rect -35 614 35 1046
rect -35 -1046 35 -614
<< ppolyres >>
rect -35 -614 35 614
<< locali >>
rect -165 1142 -69 1176
rect 69 1142 165 1176
rect -165 1080 -131 1142
rect 131 1080 165 1142
rect -165 -1142 -131 -1080
rect 131 -1142 165 -1080
rect -165 -1176 -69 -1142
rect 69 -1176 165 -1142
<< viali >>
rect -19 631 19 1028
rect -19 -1028 19 -631
<< metal1 >>
rect -25 1028 25 1040
rect -25 631 -19 1028
rect 19 631 25 1028
rect -25 619 25 631
rect -25 -631 25 -619
rect -25 -1028 -19 -631
rect 19 -1028 25 -631
rect -25 -1040 25 -1028
<< properties >>
string FIXED_BBOX -148 -1159 148 1159
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 6.3 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 6.869k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
