magic
tech sky130A
magscale 1 2
timestamp 1750694133
<< viali >>
rect 2973 7497 3007 7531
rect 3341 7497 3375 7531
rect 4353 7497 4387 7531
rect 5733 7497 5767 7531
rect 6837 7497 6871 7531
rect 2329 7429 2363 7463
rect 2697 7429 2731 7463
rect 4169 7429 4203 7463
rect 4721 7429 4755 7463
rect 6561 7429 6595 7463
rect 3157 7361 3191 7395
rect 3617 7361 3651 7395
rect 4537 7361 4571 7395
rect 5089 7361 5123 7395
rect 5641 7361 5675 7395
rect 6193 7361 6227 7395
rect 6745 7361 6779 7395
rect 3893 7293 3927 7327
rect 3985 6953 4019 6987
rect 5549 6953 5583 6987
rect 4261 6885 4295 6919
rect 5089 6885 5123 6919
rect 2421 6817 2455 6851
rect 3433 6749 3467 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 4905 6749 4939 6783
rect 5549 6749 5583 6783
rect 5825 6749 5859 6783
rect 7573 6749 7607 6783
rect 2697 6681 2731 6715
rect 3249 6681 3283 6715
rect 3801 6681 3835 6715
rect 5273 6681 5307 6715
rect 5457 6681 5491 6715
rect 7205 6681 7239 6715
rect 2973 6613 3007 6647
rect 5641 6613 5675 6647
rect 2329 6409 2363 6443
rect 3985 6409 4019 6443
rect 4721 6409 4755 6443
rect 5733 6409 5767 6443
rect 6285 6409 6319 6443
rect 2605 6273 2639 6307
rect 2697 6273 2731 6307
rect 2789 6273 2823 6307
rect 3433 6273 3467 6307
rect 4169 6273 4203 6307
rect 5365 6273 5399 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 5917 6273 5951 6307
rect 6009 6273 6043 6307
rect 6101 6273 6135 6307
rect 3065 6205 3099 6239
rect 3709 6205 3743 6239
rect 4445 6205 4479 6239
rect 3341 6137 3375 6171
rect 2697 6069 2731 6103
rect 2973 6069 3007 6103
rect 3801 6069 3835 6103
rect 4261 6069 4295 6103
rect 3065 5865 3099 5899
rect 3249 5865 3283 5899
rect 3893 5865 3927 5899
rect 5181 5865 5215 5899
rect 3617 5797 3651 5831
rect 4261 5661 4295 5695
rect 4813 5661 4847 5695
rect 4905 5661 4939 5695
rect 4997 5661 5031 5695
rect 2697 5593 2731 5627
rect 3249 5593 3283 5627
rect 2421 5525 2455 5559
rect 3709 5525 3743 5559
rect 3893 5525 3927 5559
rect 2605 5321 2639 5355
rect 3801 5321 3835 5355
rect 3157 5253 3191 5287
rect 3357 5253 3391 5287
rect 3617 5185 3651 5219
rect 2789 5117 2823 5151
rect 2881 5117 2915 5151
rect 2973 5117 3007 5151
rect 3525 5049 3559 5083
rect 3341 4981 3375 5015
rect 2329 4505 2363 4539
rect 2697 4505 2731 4539
rect 3525 4233 3559 4267
rect 4629 4233 4663 4267
rect 3249 4165 3283 4199
rect 2881 4097 2915 4131
rect 3709 4097 3743 4131
rect 4537 4097 4571 4131
rect 3433 3961 3467 3995
rect 3249 3893 3283 3927
rect 3985 3621 4019 3655
rect 2789 3553 2823 3587
rect 2881 3553 2915 3587
rect 4445 3553 4479 3587
rect 2973 3485 3007 3519
rect 3341 3485 3375 3519
rect 3433 3485 3467 3519
rect 3525 3485 3559 3519
rect 3801 3417 3835 3451
rect 4261 3417 4295 3451
rect 2605 3349 2639 3383
rect 3157 3349 3191 3383
rect 2329 3077 2363 3111
rect 2697 3077 2731 3111
rect 3157 3077 3191 3111
rect 2881 3009 2915 3043
rect 2973 2873 3007 2907
rect 3065 2805 3099 2839
rect 3617 2601 3651 2635
rect 5089 2601 5123 2635
rect 7389 2601 7423 2635
rect 2973 2397 3007 2431
rect 3433 2397 3467 2431
rect 5273 2397 5307 2431
rect 7573 2397 7607 2431
rect 2329 2329 2363 2363
rect 2697 2329 2731 2363
rect 3065 2261 3099 2295
<< metal1 >>
rect 2024 7642 8072 7664
rect 2024 7590 3342 7642
rect 3394 7590 3406 7642
rect 3458 7590 3470 7642
rect 3522 7590 3534 7642
rect 3586 7590 3598 7642
rect 3650 7590 4814 7642
rect 4866 7590 4878 7642
rect 4930 7590 4942 7642
rect 4994 7590 5006 7642
rect 5058 7590 5070 7642
rect 5122 7590 6286 7642
rect 6338 7590 6350 7642
rect 6402 7590 6414 7642
rect 6466 7590 6478 7642
rect 6530 7590 6542 7642
rect 6594 7590 7758 7642
rect 7810 7590 7822 7642
rect 7874 7590 7886 7642
rect 7938 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8072 7642
rect 2024 7568 8072 7590
rect 2961 7531 3019 7537
rect 2961 7497 2973 7531
rect 3007 7497 3019 7531
rect 2961 7491 3019 7497
rect 842 7420 848 7472
rect 900 7460 906 7472
rect 2317 7463 2375 7469
rect 2317 7460 2329 7463
rect 900 7432 2329 7460
rect 900 7420 906 7432
rect 2317 7429 2329 7432
rect 2363 7429 2375 7463
rect 2317 7423 2375 7429
rect 2685 7463 2743 7469
rect 2685 7429 2697 7463
rect 2731 7460 2743 7463
rect 2976 7460 3004 7491
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 3200 7500 3341 7528
rect 3200 7488 3206 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 3329 7491 3387 7497
rect 4172 7500 4353 7528
rect 4172 7469 4200 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5592 7500 5733 7528
rect 5592 7488 5598 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 2731 7432 3004 7460
rect 4157 7463 4215 7469
rect 2731 7429 2743 7432
rect 2685 7423 2743 7429
rect 4157 7429 4169 7463
rect 4203 7429 4215 7463
rect 4157 7423 4215 7429
rect 4614 7420 4620 7472
rect 4672 7460 4678 7472
rect 4709 7463 4767 7469
rect 4709 7460 4721 7463
rect 4672 7432 4721 7460
rect 4672 7420 4678 7432
rect 4709 7429 4721 7432
rect 4755 7429 4767 7463
rect 4709 7423 4767 7429
rect 6549 7463 6607 7469
rect 6549 7429 6561 7463
rect 6595 7460 6607 7463
rect 9122 7460 9128 7472
rect 6595 7432 9128 7460
rect 6595 7429 6607 7432
rect 6549 7423 6607 7429
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5166 7392 5172 7404
rect 5123 7364 5172 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 5902 7392 5908 7404
rect 5675 7364 5908 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 2004 7296 3893 7324
rect 2004 7284 2010 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 2024 7098 7912 7120
rect 2024 7046 2606 7098
rect 2658 7046 2670 7098
rect 2722 7046 2734 7098
rect 2786 7046 2798 7098
rect 2850 7046 2862 7098
rect 2914 7046 4078 7098
rect 4130 7046 4142 7098
rect 4194 7046 4206 7098
rect 4258 7046 4270 7098
rect 4322 7046 4334 7098
rect 4386 7046 5550 7098
rect 5602 7046 5614 7098
rect 5666 7046 5678 7098
rect 5730 7046 5742 7098
rect 5794 7046 5806 7098
rect 5858 7046 7022 7098
rect 7074 7046 7086 7098
rect 7138 7046 7150 7098
rect 7202 7046 7214 7098
rect 7266 7046 7278 7098
rect 7330 7046 7912 7098
rect 2024 7024 7912 7046
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 3973 6987 4031 6993
rect 3973 6984 3985 6987
rect 3660 6956 3985 6984
rect 3660 6944 3666 6956
rect 3973 6953 3985 6956
rect 4019 6953 4031 6987
rect 3973 6947 4031 6953
rect 5537 6987 5595 6993
rect 5537 6953 5549 6987
rect 5583 6984 5595 6987
rect 6178 6984 6184 6996
rect 5583 6956 6184 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 4249 6919 4307 6925
rect 4249 6885 4261 6919
rect 4295 6885 4307 6919
rect 4249 6879 4307 6885
rect 5077 6919 5135 6925
rect 5077 6885 5089 6919
rect 5123 6885 5135 6919
rect 5077 6879 5135 6885
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2958 6848 2964 6860
rect 2455 6820 2964 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 4264 6848 4292 6879
rect 3528 6820 4292 6848
rect 5092 6848 5120 6879
rect 5902 6848 5908 6860
rect 5092 6820 5908 6848
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 1360 6752 3433 6780
rect 1360 6740 1366 6752
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 2685 6715 2743 6721
rect 2685 6681 2697 6715
rect 2731 6712 2743 6715
rect 3237 6715 3295 6721
rect 2731 6684 3188 6712
rect 2731 6681 2743 6684
rect 2685 6675 2743 6681
rect 750 6604 756 6656
rect 808 6644 814 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 808 6616 2973 6644
rect 808 6604 814 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 3160 6644 3188 6684
rect 3237 6681 3249 6715
rect 3283 6712 3295 6715
rect 3528 6712 3556 6820
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 4028 6752 4169 6780
rect 4028 6740 4034 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4430 6740 4436 6792
rect 4488 6740 4494 6792
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4764 6752 4905 6780
rect 4764 6740 4770 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 3283 6684 3556 6712
rect 3283 6681 3295 6684
rect 3237 6675 3295 6681
rect 3786 6672 3792 6724
rect 3844 6672 3850 6724
rect 5258 6672 5264 6724
rect 5316 6672 5322 6724
rect 5442 6672 5448 6724
rect 5500 6672 5506 6724
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 7193 6715 7251 6721
rect 7193 6712 7205 6715
rect 5776 6684 7205 6712
rect 5776 6672 5782 6684
rect 7193 6681 7205 6684
rect 7239 6681 7251 6715
rect 7193 6675 7251 6681
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 3160 6616 5641 6644
rect 2961 6607 3019 6613
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 2024 6554 8072 6576
rect 2024 6502 3342 6554
rect 3394 6502 3406 6554
rect 3458 6502 3470 6554
rect 3522 6502 3534 6554
rect 3586 6502 3598 6554
rect 3650 6502 4814 6554
rect 4866 6502 4878 6554
rect 4930 6502 4942 6554
rect 4994 6502 5006 6554
rect 5058 6502 5070 6554
rect 5122 6502 6286 6554
rect 6338 6502 6350 6554
rect 6402 6502 6414 6554
rect 6466 6502 6478 6554
rect 6530 6502 6542 6554
rect 6594 6502 7758 6554
rect 7810 6502 7822 6554
rect 7874 6502 7886 6554
rect 7938 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8072 6554
rect 2024 6480 8072 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6409 2375 6443
rect 2317 6403 2375 6409
rect 2332 6372 2360 6403
rect 2590 6400 2596 6452
rect 2648 6440 2654 6452
rect 3050 6440 3056 6452
rect 2648 6412 3056 6440
rect 2648 6400 2654 6412
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 3970 6400 3976 6452
rect 4028 6400 4034 6452
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 5442 6440 5448 6452
rect 5368 6412 5448 6440
rect 4430 6372 4436 6384
rect 2332 6344 4436 6372
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 2590 6264 2596 6316
rect 2648 6264 2654 6316
rect 2682 6264 2688 6316
rect 2740 6264 2746 6316
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 2823 6276 2912 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2884 6168 2912 6276
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3234 6304 3240 6316
rect 3016 6276 3240 6304
rect 3016 6264 3022 6276
rect 3234 6264 3240 6276
rect 3292 6304 3298 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3292 6276 3433 6304
rect 3292 6264 3298 6276
rect 3421 6273 3433 6276
rect 3467 6304 3479 6307
rect 4062 6304 4068 6316
rect 3467 6276 4068 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4614 6304 4620 6316
rect 4203 6276 4620 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5368 6313 5396 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 5718 6400 5724 6452
rect 5776 6400 5782 6452
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 6730 6440 6736 6452
rect 6319 6412 6736 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 5552 6372 5580 6400
rect 5460 6344 6040 6372
rect 5460 6316 5488 6344
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 3050 6196 3056 6248
rect 3108 6236 3114 6248
rect 3602 6236 3608 6248
rect 3108 6208 3608 6236
rect 3108 6196 3114 6208
rect 3602 6196 3608 6208
rect 3660 6236 3666 6248
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3660 6208 3709 6236
rect 3660 6196 3666 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 3936 6208 4445 6236
rect 3936 6196 3942 6208
rect 4433 6205 4445 6208
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 3329 6171 3387 6177
rect 2700 6140 3096 6168
rect 2700 6109 2728 6140
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6069 2743 6103
rect 2685 6063 2743 6069
rect 2958 6060 2964 6112
rect 3016 6060 3022 6112
rect 3068 6100 3096 6140
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 4522 6168 4528 6180
rect 3375 6140 4528 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 4982 6128 4988 6180
rect 5040 6168 5046 6180
rect 5368 6168 5396 6267
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6012 6313 6040 6344
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 5592 6276 5917 6304
rect 5592 6264 5598 6276
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6104 6168 6132 6267
rect 5040 6140 6132 6168
rect 5040 6128 5046 6140
rect 3789 6103 3847 6109
rect 3789 6100 3801 6103
rect 3068 6072 3801 6100
rect 3789 6069 3801 6072
rect 3835 6100 3847 6103
rect 3878 6100 3884 6112
rect 3835 6072 3884 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 4120 6072 4261 6100
rect 4120 6060 4126 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 5258 6060 5264 6112
rect 5316 6100 5322 6112
rect 5442 6100 5448 6112
rect 5316 6072 5448 6100
rect 5316 6060 5322 6072
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 2024 6010 7912 6032
rect 2024 5958 2606 6010
rect 2658 5958 2670 6010
rect 2722 5958 2734 6010
rect 2786 5958 2798 6010
rect 2850 5958 2862 6010
rect 2914 5958 4078 6010
rect 4130 5958 4142 6010
rect 4194 5958 4206 6010
rect 4258 5958 4270 6010
rect 4322 5958 4334 6010
rect 4386 5958 5550 6010
rect 5602 5958 5614 6010
rect 5666 5958 5678 6010
rect 5730 5958 5742 6010
rect 5794 5958 5806 6010
rect 5858 5958 7022 6010
rect 7074 5958 7086 6010
rect 7138 5958 7150 6010
rect 7202 5958 7214 6010
rect 7266 5958 7278 6010
rect 7330 5958 7912 6010
rect 2024 5936 7912 5958
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3142 5896 3148 5908
rect 3099 5868 3148 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 3878 5856 3884 5908
rect 3936 5856 3942 5908
rect 5166 5856 5172 5908
rect 5224 5856 5230 5908
rect 3605 5831 3663 5837
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 3970 5828 3976 5840
rect 3651 5800 3976 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 3970 5788 3976 5800
rect 4028 5828 4034 5840
rect 4982 5828 4988 5840
rect 4028 5800 4988 5828
rect 4028 5788 4034 5800
rect 4982 5788 4988 5800
rect 5040 5788 5046 5840
rect 5350 5760 5356 5772
rect 4816 5732 5356 5760
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4120 5664 4261 5692
rect 4120 5652 4126 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 2682 5584 2688 5636
rect 2740 5584 2746 5636
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 3602 5624 3608 5636
rect 3283 5596 3608 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 3602 5584 3608 5596
rect 3660 5624 3666 5636
rect 4264 5624 4292 5655
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 4816 5701 4844 5732
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4764 5664 4813 5692
rect 4764 5652 4770 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 4908 5624 4936 5655
rect 4982 5652 4988 5704
rect 5040 5652 5046 5704
rect 5442 5624 5448 5636
rect 3660 5596 3924 5624
rect 4264 5596 5448 5624
rect 3660 5584 3666 5596
rect 2406 5516 2412 5568
rect 2464 5516 2470 5568
rect 3694 5516 3700 5568
rect 3752 5516 3758 5568
rect 3896 5565 3924 5596
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 4522 5556 4528 5568
rect 3927 5528 4528 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 2024 5466 8072 5488
rect 2024 5414 3342 5466
rect 3394 5414 3406 5466
rect 3458 5414 3470 5466
rect 3522 5414 3534 5466
rect 3586 5414 3598 5466
rect 3650 5414 4814 5466
rect 4866 5414 4878 5466
rect 4930 5414 4942 5466
rect 4994 5414 5006 5466
rect 5058 5414 5070 5466
rect 5122 5414 6286 5466
rect 6338 5414 6350 5466
rect 6402 5414 6414 5466
rect 6466 5414 6478 5466
rect 6530 5414 6542 5466
rect 6594 5414 7758 5466
rect 7810 5414 7822 5466
rect 7874 5414 7886 5466
rect 7938 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8072 5466
rect 2024 5392 8072 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 2682 5352 2688 5364
rect 2639 5324 2688 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 2792 5324 3372 5352
rect 2792 5157 2820 5324
rect 3344 5293 3372 5324
rect 3786 5312 3792 5364
rect 3844 5312 3850 5364
rect 3145 5287 3203 5293
rect 3145 5253 3157 5287
rect 3191 5253 3203 5287
rect 3344 5287 3403 5293
rect 3344 5256 3357 5287
rect 3145 5247 3203 5253
rect 3345 5253 3357 5256
rect 3391 5284 3403 5287
rect 4062 5284 4068 5296
rect 3391 5256 4068 5284
rect 3391 5253 3403 5256
rect 3345 5247 3403 5253
rect 3160 5160 3188 5247
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3694 5216 3700 5228
rect 3651 5188 3700 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5117 2835 5151
rect 2777 5111 2835 5117
rect 2792 5080 2820 5111
rect 2866 5108 2872 5160
rect 2924 5108 2930 5160
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3142 5148 3148 5160
rect 3007 5120 3148 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3142 5108 3148 5120
rect 3200 5148 3206 5160
rect 4706 5148 4712 5160
rect 3200 5120 4712 5148
rect 3200 5108 3206 5120
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 3513 5083 3571 5089
rect 2792 5052 3004 5080
rect 2976 5024 3004 5052
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 5902 5080 5908 5092
rect 3559 5052 5908 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 2958 4972 2964 5024
rect 3016 4972 3022 5024
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 3329 5015 3387 5021
rect 3329 5012 3341 5015
rect 3108 4984 3341 5012
rect 3108 4972 3114 4984
rect 3329 4981 3341 4984
rect 3375 5012 3387 5015
rect 3970 5012 3976 5024
rect 3375 4984 3976 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 2024 4922 7912 4944
rect 2024 4870 2606 4922
rect 2658 4870 2670 4922
rect 2722 4870 2734 4922
rect 2786 4870 2798 4922
rect 2850 4870 2862 4922
rect 2914 4870 4078 4922
rect 4130 4870 4142 4922
rect 4194 4870 4206 4922
rect 4258 4870 4270 4922
rect 4322 4870 4334 4922
rect 4386 4870 5550 4922
rect 5602 4870 5614 4922
rect 5666 4870 5678 4922
rect 5730 4870 5742 4922
rect 5794 4870 5806 4922
rect 5858 4870 7022 4922
rect 7074 4870 7086 4922
rect 7138 4870 7150 4922
rect 7202 4870 7214 4922
rect 7266 4870 7278 4922
rect 7330 4870 7912 4922
rect 2024 4848 7912 4870
rect 1210 4496 1216 4548
rect 1268 4536 1274 4548
rect 2317 4539 2375 4545
rect 2317 4536 2329 4539
rect 1268 4508 2329 4536
rect 1268 4496 1274 4508
rect 2317 4505 2329 4508
rect 2363 4505 2375 4539
rect 2317 4499 2375 4505
rect 2685 4539 2743 4545
rect 2685 4505 2697 4539
rect 2731 4536 2743 4539
rect 3142 4536 3148 4548
rect 2731 4508 3148 4536
rect 2731 4505 2743 4508
rect 2685 4499 2743 4505
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 2024 4378 8072 4400
rect 2024 4326 3342 4378
rect 3394 4326 3406 4378
rect 3458 4326 3470 4378
rect 3522 4326 3534 4378
rect 3586 4326 3598 4378
rect 3650 4326 4814 4378
rect 4866 4326 4878 4378
rect 4930 4326 4942 4378
rect 4994 4326 5006 4378
rect 5058 4326 5070 4378
rect 5122 4326 6286 4378
rect 6338 4326 6350 4378
rect 6402 4326 6414 4378
rect 6466 4326 6478 4378
rect 6530 4326 6542 4378
rect 6594 4326 7758 4378
rect 7810 4326 7822 4378
rect 7874 4326 7886 4378
rect 7938 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8072 4378
rect 2024 4304 8072 4326
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 3513 4267 3571 4273
rect 3513 4264 3525 4267
rect 3200 4236 3525 4264
rect 3200 4224 3206 4236
rect 3513 4233 3525 4236
rect 3559 4233 3571 4267
rect 3513 4227 3571 4233
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 4706 4264 4712 4276
rect 4663 4236 4712 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 3234 4156 3240 4208
rect 3292 4196 3298 4208
rect 4430 4196 4436 4208
rect 3292 4168 4436 4196
rect 3292 4156 3298 4168
rect 4430 4156 4436 4168
rect 4488 4156 4494 4208
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3050 4128 3056 4140
rect 2915 4100 3056 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3436 4100 3709 4128
rect 3436 4001 3464 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 7374 4128 7380 4140
rect 4580 4100 7380 4128
rect 4580 4088 4586 4100
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 3421 3995 3479 4001
rect 3421 3961 3433 3995
rect 3467 3961 3479 3995
rect 3421 3955 3479 3961
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3786 3924 3792 3936
rect 3283 3896 3792 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 2024 3834 7912 3856
rect 2024 3782 2606 3834
rect 2658 3782 2670 3834
rect 2722 3782 2734 3834
rect 2786 3782 2798 3834
rect 2850 3782 2862 3834
rect 2914 3782 4078 3834
rect 4130 3782 4142 3834
rect 4194 3782 4206 3834
rect 4258 3782 4270 3834
rect 4322 3782 4334 3834
rect 4386 3782 5550 3834
rect 5602 3782 5614 3834
rect 5666 3782 5678 3834
rect 5730 3782 5742 3834
rect 5794 3782 5806 3834
rect 5858 3782 7022 3834
rect 7074 3782 7086 3834
rect 7138 3782 7150 3834
rect 7202 3782 7214 3834
rect 7266 3782 7278 3834
rect 7330 3782 7912 3834
rect 2024 3760 7912 3782
rect 3970 3652 3976 3664
rect 2792 3624 3976 3652
rect 2792 3596 2820 3624
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 2774 3544 2780 3596
rect 2832 3544 2838 3596
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 3050 3584 3056 3596
rect 2915 3556 3056 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 3344 3556 4445 3584
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3344 3525 3372 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3016 3488 3341 3516
rect 3016 3476 3022 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3970 3516 3976 3528
rect 3559 3488 3976 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 3436 3448 3464 3479
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 3108 3420 3464 3448
rect 3108 3408 3114 3420
rect 3786 3408 3792 3460
rect 3844 3408 3850 3460
rect 4249 3451 4307 3457
rect 4249 3417 4261 3451
rect 4295 3448 4307 3451
rect 4430 3448 4436 3460
rect 4295 3420 4436 3448
rect 4295 3417 4307 3420
rect 4249 3411 4307 3417
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 2593 3383 2651 3389
rect 2593 3349 2605 3383
rect 2639 3380 2651 3383
rect 2682 3380 2688 3392
rect 2639 3352 2688 3380
rect 2639 3349 2651 3352
rect 2593 3343 2651 3349
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 3142 3340 3148 3392
rect 3200 3340 3206 3392
rect 2024 3290 8072 3312
rect 2024 3238 3342 3290
rect 3394 3238 3406 3290
rect 3458 3238 3470 3290
rect 3522 3238 3534 3290
rect 3586 3238 3598 3290
rect 3650 3238 4814 3290
rect 4866 3238 4878 3290
rect 4930 3238 4942 3290
rect 4994 3238 5006 3290
rect 5058 3238 5070 3290
rect 5122 3238 6286 3290
rect 6338 3238 6350 3290
rect 6402 3238 6414 3290
rect 6466 3238 6478 3290
rect 6530 3238 6542 3290
rect 6594 3238 7758 3290
rect 7810 3238 7822 3290
rect 7874 3238 7886 3290
rect 7938 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8072 3290
rect 2024 3216 8072 3238
rect 1210 3068 1216 3120
rect 1268 3108 1274 3120
rect 2317 3111 2375 3117
rect 2317 3108 2329 3111
rect 1268 3080 2329 3108
rect 1268 3068 1274 3080
rect 2317 3077 2329 3080
rect 2363 3077 2375 3111
rect 2317 3071 2375 3077
rect 2682 3068 2688 3120
rect 2740 3068 2746 3120
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 3145 3111 3203 3117
rect 3145 3108 3157 3111
rect 3108 3080 3157 3108
rect 3108 3068 3114 3080
rect 3145 3077 3157 3080
rect 3191 3077 3203 3111
rect 3145 3071 3203 3077
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 2958 3040 2964 3052
rect 2915 3012 2964 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 2774 2864 2780 2916
rect 2832 2904 2838 2916
rect 2961 2907 3019 2913
rect 2961 2904 2973 2907
rect 2832 2876 2973 2904
rect 2832 2864 2838 2876
rect 2961 2873 2973 2876
rect 3007 2873 3019 2907
rect 2961 2867 3019 2873
rect 3050 2796 3056 2848
rect 3108 2796 3114 2848
rect 2024 2746 7912 2768
rect 2024 2694 2606 2746
rect 2658 2694 2670 2746
rect 2722 2694 2734 2746
rect 2786 2694 2798 2746
rect 2850 2694 2862 2746
rect 2914 2694 4078 2746
rect 4130 2694 4142 2746
rect 4194 2694 4206 2746
rect 4258 2694 4270 2746
rect 4322 2694 4334 2746
rect 4386 2694 5550 2746
rect 5602 2694 5614 2746
rect 5666 2694 5678 2746
rect 5730 2694 5742 2746
rect 5794 2694 5806 2746
rect 5858 2694 7022 2746
rect 7074 2694 7086 2746
rect 7138 2694 7150 2746
rect 7202 2694 7214 2746
rect 7266 2694 7278 2746
rect 7330 2694 7912 2746
rect 2024 2672 7912 2694
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3786 2632 3792 2644
rect 3651 2604 3792 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4430 2592 4436 2644
rect 4488 2632 4494 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4488 2604 5089 2632
rect 4488 2592 4494 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 1670 2456 1676 2508
rect 1728 2496 1734 2508
rect 1728 2468 3464 2496
rect 1728 2456 1734 2468
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3050 2428 3056 2440
rect 3007 2400 3056 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3436 2437 3464 2468
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 5224 2400 5273 2428
rect 5224 2388 5230 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8294 2428 8300 2440
rect 7607 2400 8300 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2317 2363 2375 2369
rect 2317 2360 2329 2363
rect 1268 2332 2329 2360
rect 1268 2320 1274 2332
rect 2317 2329 2329 2332
rect 2363 2329 2375 2363
rect 2317 2323 2375 2329
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 3142 2360 3148 2372
rect 2731 2332 3148 2360
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 3142 2320 3148 2332
rect 3200 2320 3206 2372
rect 3050 2252 3056 2304
rect 3108 2252 3114 2304
rect 2024 2202 8072 2224
rect 2024 2150 3342 2202
rect 3394 2150 3406 2202
rect 3458 2150 3470 2202
rect 3522 2150 3534 2202
rect 3586 2150 3598 2202
rect 3650 2150 4814 2202
rect 4866 2150 4878 2202
rect 4930 2150 4942 2202
rect 4994 2150 5006 2202
rect 5058 2150 5070 2202
rect 5122 2150 6286 2202
rect 6338 2150 6350 2202
rect 6402 2150 6414 2202
rect 6466 2150 6478 2202
rect 6530 2150 6542 2202
rect 6594 2150 7758 2202
rect 7810 2150 7822 2202
rect 7874 2150 7886 2202
rect 7938 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8072 2202
rect 2024 2128 8072 2150
<< via1 >>
rect 3342 7590 3394 7642
rect 3406 7590 3458 7642
rect 3470 7590 3522 7642
rect 3534 7590 3586 7642
rect 3598 7590 3650 7642
rect 4814 7590 4866 7642
rect 4878 7590 4930 7642
rect 4942 7590 4994 7642
rect 5006 7590 5058 7642
rect 5070 7590 5122 7642
rect 6286 7590 6338 7642
rect 6350 7590 6402 7642
rect 6414 7590 6466 7642
rect 6478 7590 6530 7642
rect 6542 7590 6594 7642
rect 7758 7590 7810 7642
rect 7822 7590 7874 7642
rect 7886 7590 7938 7642
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 848 7420 900 7472
rect 3148 7488 3200 7540
rect 5540 7488 5592 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 4620 7420 4672 7472
rect 9128 7420 9180 7472
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 5172 7352 5224 7404
rect 5908 7352 5960 7404
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 1952 7284 2004 7336
rect 2606 7046 2658 7098
rect 2670 7046 2722 7098
rect 2734 7046 2786 7098
rect 2798 7046 2850 7098
rect 2862 7046 2914 7098
rect 4078 7046 4130 7098
rect 4142 7046 4194 7098
rect 4206 7046 4258 7098
rect 4270 7046 4322 7098
rect 4334 7046 4386 7098
rect 5550 7046 5602 7098
rect 5614 7046 5666 7098
rect 5678 7046 5730 7098
rect 5742 7046 5794 7098
rect 5806 7046 5858 7098
rect 7022 7046 7074 7098
rect 7086 7046 7138 7098
rect 7150 7046 7202 7098
rect 7214 7046 7266 7098
rect 7278 7046 7330 7098
rect 3608 6944 3660 6996
rect 6184 6944 6236 6996
rect 2964 6808 3016 6860
rect 1308 6740 1360 6792
rect 756 6604 808 6656
rect 5908 6808 5960 6860
rect 3976 6740 4028 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4712 6740 4764 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 3792 6715 3844 6724
rect 3792 6681 3801 6715
rect 3801 6681 3835 6715
rect 3835 6681 3844 6715
rect 3792 6672 3844 6681
rect 5264 6715 5316 6724
rect 5264 6681 5273 6715
rect 5273 6681 5307 6715
rect 5307 6681 5316 6715
rect 5264 6672 5316 6681
rect 5448 6715 5500 6724
rect 5448 6681 5457 6715
rect 5457 6681 5491 6715
rect 5491 6681 5500 6715
rect 5448 6672 5500 6681
rect 5724 6672 5776 6724
rect 3342 6502 3394 6554
rect 3406 6502 3458 6554
rect 3470 6502 3522 6554
rect 3534 6502 3586 6554
rect 3598 6502 3650 6554
rect 4814 6502 4866 6554
rect 4878 6502 4930 6554
rect 4942 6502 4994 6554
rect 5006 6502 5058 6554
rect 5070 6502 5122 6554
rect 6286 6502 6338 6554
rect 6350 6502 6402 6554
rect 6414 6502 6466 6554
rect 6478 6502 6530 6554
rect 6542 6502 6594 6554
rect 7758 6502 7810 6554
rect 7822 6502 7874 6554
rect 7886 6502 7938 6554
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 2596 6400 2648 6452
rect 3056 6400 3108 6452
rect 3976 6443 4028 6452
rect 3976 6409 3985 6443
rect 3985 6409 4019 6443
rect 4019 6409 4028 6443
rect 3976 6400 4028 6409
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 4436 6332 4488 6384
rect 2596 6307 2648 6316
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 2964 6264 3016 6316
rect 3240 6264 3292 6316
rect 4068 6264 4120 6316
rect 4620 6264 4672 6316
rect 5448 6400 5500 6452
rect 5540 6400 5592 6452
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 6736 6400 6788 6452
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 3608 6196 3660 6248
rect 3884 6196 3936 6248
rect 2964 6103 3016 6112
rect 2964 6069 2973 6103
rect 2973 6069 3007 6103
rect 3007 6069 3016 6103
rect 2964 6060 3016 6069
rect 4528 6128 4580 6180
rect 4988 6128 5040 6180
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 3884 6060 3936 6112
rect 4068 6060 4120 6112
rect 5264 6060 5316 6112
rect 5448 6060 5500 6112
rect 2606 5958 2658 6010
rect 2670 5958 2722 6010
rect 2734 5958 2786 6010
rect 2798 5958 2850 6010
rect 2862 5958 2914 6010
rect 4078 5958 4130 6010
rect 4142 5958 4194 6010
rect 4206 5958 4258 6010
rect 4270 5958 4322 6010
rect 4334 5958 4386 6010
rect 5550 5958 5602 6010
rect 5614 5958 5666 6010
rect 5678 5958 5730 6010
rect 5742 5958 5794 6010
rect 5806 5958 5858 6010
rect 7022 5958 7074 6010
rect 7086 5958 7138 6010
rect 7150 5958 7202 6010
rect 7214 5958 7266 6010
rect 7278 5958 7330 6010
rect 3148 5856 3200 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 3884 5899 3936 5908
rect 3884 5865 3893 5899
rect 3893 5865 3927 5899
rect 3927 5865 3936 5899
rect 3884 5856 3936 5865
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 3976 5788 4028 5840
rect 4988 5788 5040 5840
rect 4068 5652 4120 5704
rect 2688 5627 2740 5636
rect 2688 5593 2697 5627
rect 2697 5593 2731 5627
rect 2731 5593 2740 5627
rect 2688 5584 2740 5593
rect 3608 5584 3660 5636
rect 4712 5652 4764 5704
rect 5356 5720 5408 5772
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 4988 5652 5040 5661
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 3700 5559 3752 5568
rect 3700 5525 3709 5559
rect 3709 5525 3743 5559
rect 3743 5525 3752 5559
rect 3700 5516 3752 5525
rect 5448 5584 5500 5636
rect 4528 5516 4580 5568
rect 3342 5414 3394 5466
rect 3406 5414 3458 5466
rect 3470 5414 3522 5466
rect 3534 5414 3586 5466
rect 3598 5414 3650 5466
rect 4814 5414 4866 5466
rect 4878 5414 4930 5466
rect 4942 5414 4994 5466
rect 5006 5414 5058 5466
rect 5070 5414 5122 5466
rect 6286 5414 6338 5466
rect 6350 5414 6402 5466
rect 6414 5414 6466 5466
rect 6478 5414 6530 5466
rect 6542 5414 6594 5466
rect 7758 5414 7810 5466
rect 7822 5414 7874 5466
rect 7886 5414 7938 5466
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 2688 5312 2740 5364
rect 3792 5355 3844 5364
rect 3792 5321 3801 5355
rect 3801 5321 3835 5355
rect 3835 5321 3844 5355
rect 3792 5312 3844 5321
rect 4068 5244 4120 5296
rect 3700 5176 3752 5228
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 3148 5108 3200 5160
rect 4712 5108 4764 5160
rect 5908 5040 5960 5092
rect 2964 4972 3016 5024
rect 3056 4972 3108 5024
rect 3976 4972 4028 5024
rect 2606 4870 2658 4922
rect 2670 4870 2722 4922
rect 2734 4870 2786 4922
rect 2798 4870 2850 4922
rect 2862 4870 2914 4922
rect 4078 4870 4130 4922
rect 4142 4870 4194 4922
rect 4206 4870 4258 4922
rect 4270 4870 4322 4922
rect 4334 4870 4386 4922
rect 5550 4870 5602 4922
rect 5614 4870 5666 4922
rect 5678 4870 5730 4922
rect 5742 4870 5794 4922
rect 5806 4870 5858 4922
rect 7022 4870 7074 4922
rect 7086 4870 7138 4922
rect 7150 4870 7202 4922
rect 7214 4870 7266 4922
rect 7278 4870 7330 4922
rect 1216 4496 1268 4548
rect 3148 4496 3200 4548
rect 3342 4326 3394 4378
rect 3406 4326 3458 4378
rect 3470 4326 3522 4378
rect 3534 4326 3586 4378
rect 3598 4326 3650 4378
rect 4814 4326 4866 4378
rect 4878 4326 4930 4378
rect 4942 4326 4994 4378
rect 5006 4326 5058 4378
rect 5070 4326 5122 4378
rect 6286 4326 6338 4378
rect 6350 4326 6402 4378
rect 6414 4326 6466 4378
rect 6478 4326 6530 4378
rect 6542 4326 6594 4378
rect 7758 4326 7810 4378
rect 7822 4326 7874 4378
rect 7886 4326 7938 4378
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 3148 4224 3200 4276
rect 4712 4224 4764 4276
rect 3240 4199 3292 4208
rect 3240 4165 3249 4199
rect 3249 4165 3283 4199
rect 3283 4165 3292 4199
rect 3240 4156 3292 4165
rect 4436 4156 4488 4208
rect 3056 4088 3108 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 7380 4088 7432 4140
rect 3792 3884 3844 3936
rect 2606 3782 2658 3834
rect 2670 3782 2722 3834
rect 2734 3782 2786 3834
rect 2798 3782 2850 3834
rect 2862 3782 2914 3834
rect 4078 3782 4130 3834
rect 4142 3782 4194 3834
rect 4206 3782 4258 3834
rect 4270 3782 4322 3834
rect 4334 3782 4386 3834
rect 5550 3782 5602 3834
rect 5614 3782 5666 3834
rect 5678 3782 5730 3834
rect 5742 3782 5794 3834
rect 5806 3782 5858 3834
rect 7022 3782 7074 3834
rect 7086 3782 7138 3834
rect 7150 3782 7202 3834
rect 7214 3782 7266 3834
rect 7278 3782 7330 3834
rect 3976 3655 4028 3664
rect 3976 3621 3985 3655
rect 3985 3621 4019 3655
rect 4019 3621 4028 3655
rect 3976 3612 4028 3621
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 3056 3544 3108 3596
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 3056 3408 3108 3460
rect 3976 3476 4028 3528
rect 3792 3451 3844 3460
rect 3792 3417 3801 3451
rect 3801 3417 3835 3451
rect 3835 3417 3844 3451
rect 3792 3408 3844 3417
rect 4436 3408 4488 3460
rect 2688 3340 2740 3392
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 3342 3238 3394 3290
rect 3406 3238 3458 3290
rect 3470 3238 3522 3290
rect 3534 3238 3586 3290
rect 3598 3238 3650 3290
rect 4814 3238 4866 3290
rect 4878 3238 4930 3290
rect 4942 3238 4994 3290
rect 5006 3238 5058 3290
rect 5070 3238 5122 3290
rect 6286 3238 6338 3290
rect 6350 3238 6402 3290
rect 6414 3238 6466 3290
rect 6478 3238 6530 3290
rect 6542 3238 6594 3290
rect 7758 3238 7810 3290
rect 7822 3238 7874 3290
rect 7886 3238 7938 3290
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 1216 3068 1268 3120
rect 2688 3111 2740 3120
rect 2688 3077 2697 3111
rect 2697 3077 2731 3111
rect 2731 3077 2740 3111
rect 2688 3068 2740 3077
rect 3056 3068 3108 3120
rect 2964 3000 3016 3052
rect 2780 2864 2832 2916
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 2606 2694 2658 2746
rect 2670 2694 2722 2746
rect 2734 2694 2786 2746
rect 2798 2694 2850 2746
rect 2862 2694 2914 2746
rect 4078 2694 4130 2746
rect 4142 2694 4194 2746
rect 4206 2694 4258 2746
rect 4270 2694 4322 2746
rect 4334 2694 4386 2746
rect 5550 2694 5602 2746
rect 5614 2694 5666 2746
rect 5678 2694 5730 2746
rect 5742 2694 5794 2746
rect 5806 2694 5858 2746
rect 7022 2694 7074 2746
rect 7086 2694 7138 2746
rect 7150 2694 7202 2746
rect 7214 2694 7266 2746
rect 7278 2694 7330 2746
rect 3792 2592 3844 2644
rect 4436 2592 4488 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 1676 2456 1728 2508
rect 3056 2388 3108 2440
rect 5172 2388 5224 2440
rect 8300 2388 8352 2440
rect 1216 2320 1268 2372
rect 3148 2320 3200 2372
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 3342 2150 3394 2202
rect 3406 2150 3458 2202
rect 3470 2150 3522 2202
rect 3534 2150 3586 2202
rect 3598 2150 3650 2202
rect 4814 2150 4866 2202
rect 4878 2150 4930 2202
rect 4942 2150 4994 2202
rect 5006 2150 5058 2202
rect 5070 2150 5122 2202
rect 6286 2150 6338 2202
rect 6350 2150 6402 2202
rect 6414 2150 6466 2202
rect 6478 2150 6530 2202
rect 6542 2150 6594 2202
rect 7758 2150 7810 2202
rect 7822 2150 7874 2202
rect 7886 2150 7938 2202
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
<< metal2 >>
rect 754 9600 810 10000
rect 1950 9600 2006 10000
rect 3146 9600 3202 10000
rect 4342 9738 4398 10000
rect 4342 9710 4660 9738
rect 4342 9600 4398 9710
rect 768 6662 796 9600
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 860 7478 888 7647
rect 848 7472 900 7478
rect 848 7414 900 7420
rect 1964 7342 1992 9600
rect 2962 8800 3018 8809
rect 2962 8735 3018 8744
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 2606 7100 2914 7109
rect 2606 7098 2612 7100
rect 2668 7098 2692 7100
rect 2748 7098 2772 7100
rect 2828 7098 2852 7100
rect 2908 7098 2914 7100
rect 2668 7046 2670 7098
rect 2850 7046 2852 7098
rect 2606 7044 2612 7046
rect 2668 7044 2692 7046
rect 2748 7044 2772 7046
rect 2828 7044 2852 7046
rect 2908 7044 2914 7046
rect 2606 7035 2914 7044
rect 2976 6866 3004 8735
rect 3160 7546 3188 9600
rect 3342 7644 3650 7653
rect 3342 7642 3348 7644
rect 3404 7642 3428 7644
rect 3484 7642 3508 7644
rect 3564 7642 3588 7644
rect 3644 7642 3650 7644
rect 3404 7590 3406 7642
rect 3586 7590 3588 7642
rect 3342 7588 3348 7590
rect 3404 7588 3428 7590
rect 3484 7588 3508 7590
rect 3564 7588 3588 7590
rect 3644 7588 3650 7590
rect 3342 7579 3650 7588
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 4632 7478 4660 9710
rect 5538 9600 5594 10000
rect 6734 9738 6790 10000
rect 7930 9738 7986 10000
rect 6734 9710 6868 9738
rect 6734 9600 6790 9710
rect 4814 7644 5122 7653
rect 4814 7642 4820 7644
rect 4876 7642 4900 7644
rect 4956 7642 4980 7644
rect 5036 7642 5060 7644
rect 5116 7642 5122 7644
rect 4876 7590 4878 7642
rect 5058 7590 5060 7642
rect 4814 7588 4820 7590
rect 4876 7588 4900 7590
rect 4956 7588 4980 7590
rect 5036 7588 5060 7590
rect 5116 7588 5122 7590
rect 4814 7579 5122 7588
rect 5552 7546 5580 9600
rect 6286 7644 6594 7653
rect 6286 7642 6292 7644
rect 6348 7642 6372 7644
rect 6428 7642 6452 7644
rect 6508 7642 6532 7644
rect 6588 7642 6594 7644
rect 6348 7590 6350 7642
rect 6530 7590 6532 7642
rect 6286 7588 6292 7590
rect 6348 7588 6372 7590
rect 6428 7588 6452 7590
rect 6508 7588 6532 7590
rect 6588 7588 6594 7590
rect 6286 7579 6594 7588
rect 6840 7546 6868 9710
rect 7576 9710 7986 9738
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 756 6656 808 6662
rect 1320 6633 1348 6734
rect 756 6598 808 6604
rect 1306 6624 1362 6633
rect 1306 6559 1362 6568
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2608 6322 2636 6394
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2688 6316 2740 6322
rect 2964 6316 3016 6322
rect 2740 6276 2964 6304
rect 2688 6258 2740 6264
rect 2964 6258 3016 6264
rect 2976 6118 3004 6258
rect 3068 6254 3096 6394
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2606 6012 2914 6021
rect 2606 6010 2612 6012
rect 2668 6010 2692 6012
rect 2748 6010 2772 6012
rect 2828 6010 2852 6012
rect 2908 6010 2914 6012
rect 2668 5958 2670 6010
rect 2850 5958 2852 6010
rect 2606 5956 2612 5958
rect 2668 5956 2692 5958
rect 2748 5956 2772 5958
rect 2828 5956 2852 5958
rect 2908 5956 2914 5958
rect 2606 5947 2914 5956
rect 3160 5914 3188 7346
rect 3620 7002 3648 7346
rect 4078 7100 4386 7109
rect 4078 7098 4084 7100
rect 4140 7098 4164 7100
rect 4220 7098 4244 7100
rect 4300 7098 4324 7100
rect 4380 7098 4386 7100
rect 4140 7046 4142 7098
rect 4322 7046 4324 7098
rect 4078 7044 4084 7046
rect 4140 7044 4164 7046
rect 4220 7044 4244 7046
rect 4300 7044 4324 7046
rect 4380 7044 4386 7046
rect 4078 7035 4386 7044
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3342 6556 3650 6565
rect 3342 6554 3348 6556
rect 3404 6554 3428 6556
rect 3484 6554 3508 6556
rect 3564 6554 3588 6556
rect 3644 6554 3650 6556
rect 3404 6502 3406 6554
rect 3586 6502 3588 6554
rect 3342 6500 3348 6502
rect 3404 6500 3428 6502
rect 3484 6500 3508 6502
rect 3564 6500 3588 6502
rect 3644 6500 3650 6502
rect 3342 6491 3650 6500
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3252 5914 3280 6258
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2412 5568 2464 5574
rect 2410 5536 2412 5545
rect 2464 5536 2466 5545
rect 2410 5471 2466 5480
rect 2700 5370 2728 5578
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2872 5160 2924 5166
rect 3148 5160 3200 5166
rect 2924 5108 3096 5114
rect 2872 5102 3096 5108
rect 3148 5102 3200 5108
rect 2884 5086 3096 5102
rect 3068 5030 3096 5086
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2606 4924 2914 4933
rect 2606 4922 2612 4924
rect 2668 4922 2692 4924
rect 2748 4922 2772 4924
rect 2828 4922 2852 4924
rect 2908 4922 2914 4924
rect 2668 4870 2670 4922
rect 2850 4870 2852 4922
rect 2606 4868 2612 4870
rect 2668 4868 2692 4870
rect 2748 4868 2772 4870
rect 2828 4868 2852 4870
rect 2908 4868 2914 4870
rect 2606 4859 2914 4868
rect 1216 4548 1268 4554
rect 1216 4490 1268 4496
rect 1228 4457 1256 4490
rect 1214 4448 1270 4457
rect 1214 4383 1270 4392
rect 2606 3836 2914 3845
rect 2606 3834 2612 3836
rect 2668 3834 2692 3836
rect 2748 3834 2772 3836
rect 2828 3834 2852 3836
rect 2908 3834 2914 3836
rect 2668 3782 2670 3834
rect 2850 3782 2852 3834
rect 2606 3780 2612 3782
rect 2668 3780 2692 3782
rect 2748 3780 2772 3782
rect 2828 3780 2852 3782
rect 2908 3780 2914 3782
rect 2606 3771 2914 3780
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2688 3392 2740 3398
rect 1214 3360 1270 3369
rect 2688 3334 2740 3340
rect 1214 3295 1270 3304
rect 1228 3126 1256 3295
rect 2700 3126 2728 3334
rect 1216 3120 1268 3126
rect 1216 3062 1268 3068
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2792 2922 2820 3538
rect 2976 3534 3004 4966
rect 3160 4706 3188 5102
rect 3068 4678 3188 4706
rect 3068 4146 3096 4678
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3160 4282 3188 4490
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3252 4214 3280 5850
rect 3620 5642 3648 6190
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3342 5468 3650 5477
rect 3342 5466 3348 5468
rect 3404 5466 3428 5468
rect 3484 5466 3508 5468
rect 3564 5466 3588 5468
rect 3644 5466 3650 5468
rect 3404 5414 3406 5466
rect 3586 5414 3588 5466
rect 3342 5412 3348 5414
rect 3404 5412 3428 5414
rect 3484 5412 3508 5414
rect 3564 5412 3588 5414
rect 3644 5412 3650 5414
rect 3342 5403 3650 5412
rect 3712 5234 3740 5510
rect 3804 5370 3832 6666
rect 3988 6458 4016 6734
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 4448 6390 4476 6734
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 6118 3924 6190
rect 4080 6118 4108 6258
rect 4540 6186 4568 7346
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4724 6458 4752 6734
rect 4814 6556 5122 6565
rect 4814 6554 4820 6556
rect 4876 6554 4900 6556
rect 4956 6554 4980 6556
rect 5036 6554 5060 6556
rect 5116 6554 5122 6556
rect 4876 6502 4878 6554
rect 5058 6502 5060 6554
rect 4814 6500 4820 6502
rect 4876 6500 4900 6502
rect 4956 6500 4980 6502
rect 5036 6500 5060 6502
rect 5116 6500 5122 6502
rect 4814 6491 5122 6500
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3896 5914 3924 6054
rect 4078 6012 4386 6021
rect 4078 6010 4084 6012
rect 4140 6010 4164 6012
rect 4220 6010 4244 6012
rect 4300 6010 4324 6012
rect 4380 6010 4386 6012
rect 4140 5958 4142 6010
rect 4322 5958 4324 6010
rect 4078 5956 4084 5958
rect 4140 5956 4164 5958
rect 4220 5956 4244 5958
rect 4300 5956 4324 5958
rect 4380 5956 4386 5958
rect 4078 5947 4386 5956
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3342 4380 3650 4389
rect 3342 4378 3348 4380
rect 3404 4378 3428 4380
rect 3484 4378 3508 4380
rect 3564 4378 3588 4380
rect 3644 4378 3650 4380
rect 3404 4326 3406 4378
rect 3586 4326 3588 4378
rect 3342 4324 3348 4326
rect 3404 4324 3428 4326
rect 3484 4324 3508 4326
rect 3564 4324 3588 4326
rect 3644 4324 3650 4326
rect 3342 4315 3650 4324
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3068 3602 3096 4082
rect 3792 3936 3844 3942
rect 3896 3924 3924 5850
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3988 5030 4016 5782
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5302 4108 5646
rect 4528 5568 4580 5574
rect 4632 5556 4660 6258
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 5000 5846 5028 6122
rect 5184 5914 5212 7346
rect 5550 7100 5858 7109
rect 5550 7098 5556 7100
rect 5612 7098 5636 7100
rect 5692 7098 5716 7100
rect 5772 7098 5796 7100
rect 5852 7098 5858 7100
rect 5612 7046 5614 7098
rect 5794 7046 5796 7098
rect 5550 7044 5556 7046
rect 5612 7044 5636 7046
rect 5692 7044 5716 7046
rect 5772 7044 5796 7046
rect 5852 7044 5858 7046
rect 5550 7035 5858 7044
rect 5920 6866 5948 7346
rect 6196 7002 6224 7346
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5276 6118 5304 6666
rect 5460 6458 5488 6666
rect 5552 6458 5580 6734
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5736 6458 5764 6666
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5448 6316 5500 6322
rect 5368 6276 5448 6304
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5000 5710 5028 5782
rect 5368 5778 5396 6276
rect 5448 6258 5500 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 6202 5580 6258
rect 5460 6174 5580 6202
rect 5828 6202 5856 6734
rect 6286 6556 6594 6565
rect 6286 6554 6292 6556
rect 6348 6554 6372 6556
rect 6428 6554 6452 6556
rect 6508 6554 6532 6556
rect 6588 6554 6594 6556
rect 6348 6502 6350 6554
rect 6530 6502 6532 6554
rect 6286 6500 6292 6502
rect 6348 6500 6372 6502
rect 6428 6500 6452 6502
rect 6508 6500 6532 6502
rect 6588 6500 6594 6502
rect 6286 6491 6594 6500
rect 6748 6458 6776 7346
rect 7022 7100 7330 7109
rect 7022 7098 7028 7100
rect 7084 7098 7108 7100
rect 7164 7098 7188 7100
rect 7244 7098 7268 7100
rect 7324 7098 7330 7100
rect 7084 7046 7086 7098
rect 7266 7046 7268 7098
rect 7022 7044 7028 7046
rect 7084 7044 7108 7046
rect 7164 7044 7188 7046
rect 7244 7044 7268 7046
rect 7324 7044 7330 7046
rect 7022 7035 7330 7044
rect 7576 6798 7604 9710
rect 7930 9600 7986 9710
rect 9126 9600 9182 10000
rect 7758 7644 8066 7653
rect 7758 7642 7764 7644
rect 7820 7642 7844 7644
rect 7900 7642 7924 7644
rect 7980 7642 8004 7644
rect 8060 7642 8066 7644
rect 7820 7590 7822 7642
rect 8002 7590 8004 7642
rect 7758 7588 7764 7590
rect 7820 7588 7844 7590
rect 7900 7588 7924 7590
rect 7980 7588 8004 7590
rect 8060 7588 8066 7590
rect 7758 7579 8066 7588
rect 9140 7478 9168 9600
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7758 6556 8066 6565
rect 7758 6554 7764 6556
rect 7820 6554 7844 6556
rect 7900 6554 7924 6556
rect 7980 6554 8004 6556
rect 8060 6554 8066 6556
rect 7820 6502 7822 6554
rect 8002 6502 8004 6554
rect 7758 6500 7764 6502
rect 7820 6500 7844 6502
rect 7900 6500 7924 6502
rect 7980 6500 8004 6502
rect 8060 6500 8066 6502
rect 7758 6491 8066 6500
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 5828 6174 5948 6202
rect 5460 6118 5488 6174
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4580 5528 4660 5556
rect 4528 5510 4580 5516
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3844 3896 3924 3924
rect 3792 3878 3844 3884
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2976 3058 3004 3470
rect 3068 3466 3096 3538
rect 3804 3466 3832 3878
rect 3988 3670 4016 4966
rect 4078 4924 4386 4933
rect 4078 4922 4084 4924
rect 4140 4922 4164 4924
rect 4220 4922 4244 4924
rect 4300 4922 4324 4924
rect 4380 4922 4386 4924
rect 4140 4870 4142 4922
rect 4322 4870 4324 4922
rect 4078 4868 4084 4870
rect 4140 4868 4164 4870
rect 4220 4868 4244 4870
rect 4300 4868 4324 4870
rect 4380 4868 4386 4870
rect 4078 4859 4386 4868
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4078 3836 4386 3845
rect 4078 3834 4084 3836
rect 4140 3834 4164 3836
rect 4220 3834 4244 3836
rect 4300 3834 4324 3836
rect 4380 3834 4386 3836
rect 4140 3782 4142 3834
rect 4322 3782 4324 3834
rect 4078 3780 4084 3782
rect 4140 3780 4164 3782
rect 4220 3780 4244 3782
rect 4300 3780 4324 3782
rect 4380 3780 4386 3782
rect 4078 3771 4386 3780
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3988 3534 4016 3606
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4448 3466 4476 4150
rect 4540 4146 4568 5510
rect 4724 5166 4752 5646
rect 5460 5642 5488 6054
rect 5550 6012 5858 6021
rect 5550 6010 5556 6012
rect 5612 6010 5636 6012
rect 5692 6010 5716 6012
rect 5772 6010 5796 6012
rect 5852 6010 5858 6012
rect 5612 5958 5614 6010
rect 5794 5958 5796 6010
rect 5550 5956 5556 5958
rect 5612 5956 5636 5958
rect 5692 5956 5716 5958
rect 5772 5956 5796 5958
rect 5852 5956 5858 5958
rect 5550 5947 5858 5956
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 4814 5468 5122 5477
rect 4814 5466 4820 5468
rect 4876 5466 4900 5468
rect 4956 5466 4980 5468
rect 5036 5466 5060 5468
rect 5116 5466 5122 5468
rect 4876 5414 4878 5466
rect 5058 5414 5060 5466
rect 4814 5412 4820 5414
rect 4876 5412 4900 5414
rect 4956 5412 4980 5414
rect 5036 5412 5060 5414
rect 5116 5412 5122 5414
rect 4814 5403 5122 5412
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4282 4752 5102
rect 5920 5098 5948 6174
rect 7022 6012 7330 6021
rect 7022 6010 7028 6012
rect 7084 6010 7108 6012
rect 7164 6010 7188 6012
rect 7244 6010 7268 6012
rect 7324 6010 7330 6012
rect 7084 5958 7086 6010
rect 7266 5958 7268 6010
rect 7022 5956 7028 5958
rect 7084 5956 7108 5958
rect 7164 5956 7188 5958
rect 7244 5956 7268 5958
rect 7324 5956 7330 5958
rect 7022 5947 7330 5956
rect 6286 5468 6594 5477
rect 6286 5466 6292 5468
rect 6348 5466 6372 5468
rect 6428 5466 6452 5468
rect 6508 5466 6532 5468
rect 6588 5466 6594 5468
rect 6348 5414 6350 5466
rect 6530 5414 6532 5466
rect 6286 5412 6292 5414
rect 6348 5412 6372 5414
rect 6428 5412 6452 5414
rect 6508 5412 6532 5414
rect 6588 5412 6594 5414
rect 6286 5403 6594 5412
rect 7758 5468 8066 5477
rect 7758 5466 7764 5468
rect 7820 5466 7844 5468
rect 7900 5466 7924 5468
rect 7980 5466 8004 5468
rect 8060 5466 8066 5468
rect 7820 5414 7822 5466
rect 8002 5414 8004 5466
rect 7758 5412 7764 5414
rect 7820 5412 7844 5414
rect 7900 5412 7924 5414
rect 7980 5412 8004 5414
rect 8060 5412 8066 5414
rect 7758 5403 8066 5412
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5550 4924 5858 4933
rect 5550 4922 5556 4924
rect 5612 4922 5636 4924
rect 5692 4922 5716 4924
rect 5772 4922 5796 4924
rect 5852 4922 5858 4924
rect 5612 4870 5614 4922
rect 5794 4870 5796 4922
rect 5550 4868 5556 4870
rect 5612 4868 5636 4870
rect 5692 4868 5716 4870
rect 5772 4868 5796 4870
rect 5852 4868 5858 4870
rect 5550 4859 5858 4868
rect 7022 4924 7330 4933
rect 7022 4922 7028 4924
rect 7084 4922 7108 4924
rect 7164 4922 7188 4924
rect 7244 4922 7268 4924
rect 7324 4922 7330 4924
rect 7084 4870 7086 4922
rect 7266 4870 7268 4922
rect 7022 4868 7028 4870
rect 7084 4868 7108 4870
rect 7164 4868 7188 4870
rect 7244 4868 7268 4870
rect 7324 4868 7330 4870
rect 7022 4859 7330 4868
rect 4814 4380 5122 4389
rect 4814 4378 4820 4380
rect 4876 4378 4900 4380
rect 4956 4378 4980 4380
rect 5036 4378 5060 4380
rect 5116 4378 5122 4380
rect 4876 4326 4878 4378
rect 5058 4326 5060 4378
rect 4814 4324 4820 4326
rect 4876 4324 4900 4326
rect 4956 4324 4980 4326
rect 5036 4324 5060 4326
rect 5116 4324 5122 4326
rect 4814 4315 5122 4324
rect 6286 4380 6594 4389
rect 6286 4378 6292 4380
rect 6348 4378 6372 4380
rect 6428 4378 6452 4380
rect 6508 4378 6532 4380
rect 6588 4378 6594 4380
rect 6348 4326 6350 4378
rect 6530 4326 6532 4378
rect 6286 4324 6292 4326
rect 6348 4324 6372 4326
rect 6428 4324 6452 4326
rect 6508 4324 6532 4326
rect 6588 4324 6594 4326
rect 6286 4315 6594 4324
rect 7758 4380 8066 4389
rect 7758 4378 7764 4380
rect 7820 4378 7844 4380
rect 7900 4378 7924 4380
rect 7980 4378 8004 4380
rect 8060 4378 8066 4380
rect 7820 4326 7822 4378
rect 8002 4326 8004 4378
rect 7758 4324 7764 4326
rect 7820 4324 7844 4326
rect 7900 4324 7924 4326
rect 7980 4324 8004 4326
rect 8060 4324 8066 4326
rect 7758 4315 8066 4324
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 5550 3836 5858 3845
rect 5550 3834 5556 3836
rect 5612 3834 5636 3836
rect 5692 3834 5716 3836
rect 5772 3834 5796 3836
rect 5852 3834 5858 3836
rect 5612 3782 5614 3834
rect 5794 3782 5796 3834
rect 5550 3780 5556 3782
rect 5612 3780 5636 3782
rect 5692 3780 5716 3782
rect 5772 3780 5796 3782
rect 5852 3780 5858 3782
rect 5550 3771 5858 3780
rect 7022 3836 7330 3845
rect 7022 3834 7028 3836
rect 7084 3834 7108 3836
rect 7164 3834 7188 3836
rect 7244 3834 7268 3836
rect 7324 3834 7330 3836
rect 7084 3782 7086 3834
rect 7266 3782 7268 3834
rect 7022 3780 7028 3782
rect 7084 3780 7108 3782
rect 7164 3780 7188 3782
rect 7244 3780 7268 3782
rect 7324 3780 7330 3782
rect 7022 3771 7330 3780
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 3068 3126 3096 3402
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2606 2748 2914 2757
rect 2606 2746 2612 2748
rect 2668 2746 2692 2748
rect 2748 2746 2772 2748
rect 2828 2746 2852 2748
rect 2908 2746 2914 2748
rect 2668 2694 2670 2746
rect 2850 2694 2852 2746
rect 2606 2692 2612 2694
rect 2668 2692 2692 2694
rect 2748 2692 2772 2694
rect 2828 2692 2852 2694
rect 2908 2692 2914 2694
rect 2606 2683 2914 2692
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1228 2281 1256 2314
rect 1214 2272 1270 2281
rect 1214 2207 1270 2216
rect 1688 400 1716 2450
rect 3068 2446 3096 2790
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3160 2378 3188 3334
rect 3342 3292 3650 3301
rect 3342 3290 3348 3292
rect 3404 3290 3428 3292
rect 3484 3290 3508 3292
rect 3564 3290 3588 3292
rect 3644 3290 3650 3292
rect 3404 3238 3406 3290
rect 3586 3238 3588 3290
rect 3342 3236 3348 3238
rect 3404 3236 3428 3238
rect 3484 3236 3508 3238
rect 3564 3236 3588 3238
rect 3644 3236 3650 3238
rect 3342 3227 3650 3236
rect 3804 2650 3832 3402
rect 4078 2748 4386 2757
rect 4078 2746 4084 2748
rect 4140 2746 4164 2748
rect 4220 2746 4244 2748
rect 4300 2746 4324 2748
rect 4380 2746 4386 2748
rect 4140 2694 4142 2746
rect 4322 2694 4324 2746
rect 4078 2692 4084 2694
rect 4140 2692 4164 2694
rect 4220 2692 4244 2694
rect 4300 2692 4324 2694
rect 4380 2692 4386 2694
rect 4078 2683 4386 2692
rect 4448 2650 4476 3402
rect 4814 3292 5122 3301
rect 4814 3290 4820 3292
rect 4876 3290 4900 3292
rect 4956 3290 4980 3292
rect 5036 3290 5060 3292
rect 5116 3290 5122 3292
rect 4876 3238 4878 3290
rect 5058 3238 5060 3290
rect 4814 3236 4820 3238
rect 4876 3236 4900 3238
rect 4956 3236 4980 3238
rect 5036 3236 5060 3238
rect 5116 3236 5122 3238
rect 4814 3227 5122 3236
rect 6286 3292 6594 3301
rect 6286 3290 6292 3292
rect 6348 3290 6372 3292
rect 6428 3290 6452 3292
rect 6508 3290 6532 3292
rect 6588 3290 6594 3292
rect 6348 3238 6350 3290
rect 6530 3238 6532 3290
rect 6286 3236 6292 3238
rect 6348 3236 6372 3238
rect 6428 3236 6452 3238
rect 6508 3236 6532 3238
rect 6588 3236 6594 3238
rect 6286 3227 6594 3236
rect 5550 2748 5858 2757
rect 5550 2746 5556 2748
rect 5612 2746 5636 2748
rect 5692 2746 5716 2748
rect 5772 2746 5796 2748
rect 5852 2746 5858 2748
rect 5612 2694 5614 2746
rect 5794 2694 5796 2746
rect 5550 2692 5556 2694
rect 5612 2692 5636 2694
rect 5692 2692 5716 2694
rect 5772 2692 5796 2694
rect 5852 2692 5858 2694
rect 5550 2683 5858 2692
rect 7022 2748 7330 2757
rect 7022 2746 7028 2748
rect 7084 2746 7108 2748
rect 7164 2746 7188 2748
rect 7244 2746 7268 2748
rect 7324 2746 7330 2748
rect 7084 2694 7086 2746
rect 7266 2694 7268 2746
rect 7022 2692 7028 2694
rect 7084 2692 7108 2694
rect 7164 2692 7188 2694
rect 7244 2692 7268 2694
rect 7324 2692 7330 2694
rect 7022 2683 7330 2692
rect 7392 2650 7420 4082
rect 7758 3292 8066 3301
rect 7758 3290 7764 3292
rect 7820 3290 7844 3292
rect 7900 3290 7924 3292
rect 7980 3290 8004 3292
rect 8060 3290 8066 3292
rect 7820 3238 7822 3290
rect 8002 3238 8004 3290
rect 7758 3236 7764 3238
rect 7820 3236 7844 3238
rect 7900 3236 7924 3238
rect 7980 3236 8004 3238
rect 8060 3236 8066 3238
rect 7758 3227 8066 3236
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 1193 3096 2246
rect 3342 2204 3650 2213
rect 3342 2202 3348 2204
rect 3404 2202 3428 2204
rect 3484 2202 3508 2204
rect 3564 2202 3588 2204
rect 3644 2202 3650 2204
rect 3404 2150 3406 2202
rect 3586 2150 3588 2202
rect 3342 2148 3348 2150
rect 3404 2148 3428 2150
rect 3484 2148 3508 2150
rect 3564 2148 3588 2150
rect 3644 2148 3650 2150
rect 3342 2139 3650 2148
rect 4814 2204 5122 2213
rect 4814 2202 4820 2204
rect 4876 2202 4900 2204
rect 4956 2202 4980 2204
rect 5036 2202 5060 2204
rect 5116 2202 5122 2204
rect 4876 2150 4878 2202
rect 5058 2150 5060 2202
rect 4814 2148 4820 2150
rect 4876 2148 4900 2150
rect 4956 2148 4980 2150
rect 5036 2148 5060 2150
rect 5116 2148 5122 2150
rect 4814 2139 5122 2148
rect 5184 1306 5212 2382
rect 6286 2204 6594 2213
rect 6286 2202 6292 2204
rect 6348 2202 6372 2204
rect 6428 2202 6452 2204
rect 6508 2202 6532 2204
rect 6588 2202 6594 2204
rect 6348 2150 6350 2202
rect 6530 2150 6532 2202
rect 6286 2148 6292 2150
rect 6348 2148 6372 2150
rect 6428 2148 6452 2150
rect 6508 2148 6532 2150
rect 6588 2148 6594 2150
rect 6286 2139 6594 2148
rect 7758 2204 8066 2213
rect 7758 2202 7764 2204
rect 7820 2202 7844 2204
rect 7900 2202 7924 2204
rect 7980 2202 8004 2204
rect 8060 2202 8066 2204
rect 7820 2150 7822 2202
rect 8002 2150 8004 2202
rect 7758 2148 7764 2150
rect 7820 2148 7844 2150
rect 7900 2148 7924 2150
rect 7980 2148 8004 2150
rect 8060 2148 8066 2150
rect 7758 2139 8066 2148
rect 5000 1278 5212 1306
rect 3054 1184 3110 1193
rect 3054 1119 3110 1128
rect 5000 400 5028 1278
rect 8312 400 8340 2382
rect 1674 0 1730 400
rect 4986 0 5042 400
rect 8298 0 8354 400
<< via2 >>
rect 846 7656 902 7712
rect 2962 8744 3018 8800
rect 2612 7098 2668 7100
rect 2692 7098 2748 7100
rect 2772 7098 2828 7100
rect 2852 7098 2908 7100
rect 2612 7046 2658 7098
rect 2658 7046 2668 7098
rect 2692 7046 2722 7098
rect 2722 7046 2734 7098
rect 2734 7046 2748 7098
rect 2772 7046 2786 7098
rect 2786 7046 2798 7098
rect 2798 7046 2828 7098
rect 2852 7046 2862 7098
rect 2862 7046 2908 7098
rect 2612 7044 2668 7046
rect 2692 7044 2748 7046
rect 2772 7044 2828 7046
rect 2852 7044 2908 7046
rect 3348 7642 3404 7644
rect 3428 7642 3484 7644
rect 3508 7642 3564 7644
rect 3588 7642 3644 7644
rect 3348 7590 3394 7642
rect 3394 7590 3404 7642
rect 3428 7590 3458 7642
rect 3458 7590 3470 7642
rect 3470 7590 3484 7642
rect 3508 7590 3522 7642
rect 3522 7590 3534 7642
rect 3534 7590 3564 7642
rect 3588 7590 3598 7642
rect 3598 7590 3644 7642
rect 3348 7588 3404 7590
rect 3428 7588 3484 7590
rect 3508 7588 3564 7590
rect 3588 7588 3644 7590
rect 4820 7642 4876 7644
rect 4900 7642 4956 7644
rect 4980 7642 5036 7644
rect 5060 7642 5116 7644
rect 4820 7590 4866 7642
rect 4866 7590 4876 7642
rect 4900 7590 4930 7642
rect 4930 7590 4942 7642
rect 4942 7590 4956 7642
rect 4980 7590 4994 7642
rect 4994 7590 5006 7642
rect 5006 7590 5036 7642
rect 5060 7590 5070 7642
rect 5070 7590 5116 7642
rect 4820 7588 4876 7590
rect 4900 7588 4956 7590
rect 4980 7588 5036 7590
rect 5060 7588 5116 7590
rect 6292 7642 6348 7644
rect 6372 7642 6428 7644
rect 6452 7642 6508 7644
rect 6532 7642 6588 7644
rect 6292 7590 6338 7642
rect 6338 7590 6348 7642
rect 6372 7590 6402 7642
rect 6402 7590 6414 7642
rect 6414 7590 6428 7642
rect 6452 7590 6466 7642
rect 6466 7590 6478 7642
rect 6478 7590 6508 7642
rect 6532 7590 6542 7642
rect 6542 7590 6588 7642
rect 6292 7588 6348 7590
rect 6372 7588 6428 7590
rect 6452 7588 6508 7590
rect 6532 7588 6588 7590
rect 1306 6568 1362 6624
rect 2612 6010 2668 6012
rect 2692 6010 2748 6012
rect 2772 6010 2828 6012
rect 2852 6010 2908 6012
rect 2612 5958 2658 6010
rect 2658 5958 2668 6010
rect 2692 5958 2722 6010
rect 2722 5958 2734 6010
rect 2734 5958 2748 6010
rect 2772 5958 2786 6010
rect 2786 5958 2798 6010
rect 2798 5958 2828 6010
rect 2852 5958 2862 6010
rect 2862 5958 2908 6010
rect 2612 5956 2668 5958
rect 2692 5956 2748 5958
rect 2772 5956 2828 5958
rect 2852 5956 2908 5958
rect 4084 7098 4140 7100
rect 4164 7098 4220 7100
rect 4244 7098 4300 7100
rect 4324 7098 4380 7100
rect 4084 7046 4130 7098
rect 4130 7046 4140 7098
rect 4164 7046 4194 7098
rect 4194 7046 4206 7098
rect 4206 7046 4220 7098
rect 4244 7046 4258 7098
rect 4258 7046 4270 7098
rect 4270 7046 4300 7098
rect 4324 7046 4334 7098
rect 4334 7046 4380 7098
rect 4084 7044 4140 7046
rect 4164 7044 4220 7046
rect 4244 7044 4300 7046
rect 4324 7044 4380 7046
rect 3348 6554 3404 6556
rect 3428 6554 3484 6556
rect 3508 6554 3564 6556
rect 3588 6554 3644 6556
rect 3348 6502 3394 6554
rect 3394 6502 3404 6554
rect 3428 6502 3458 6554
rect 3458 6502 3470 6554
rect 3470 6502 3484 6554
rect 3508 6502 3522 6554
rect 3522 6502 3534 6554
rect 3534 6502 3564 6554
rect 3588 6502 3598 6554
rect 3598 6502 3644 6554
rect 3348 6500 3404 6502
rect 3428 6500 3484 6502
rect 3508 6500 3564 6502
rect 3588 6500 3644 6502
rect 2410 5516 2412 5536
rect 2412 5516 2464 5536
rect 2464 5516 2466 5536
rect 2410 5480 2466 5516
rect 2612 4922 2668 4924
rect 2692 4922 2748 4924
rect 2772 4922 2828 4924
rect 2852 4922 2908 4924
rect 2612 4870 2658 4922
rect 2658 4870 2668 4922
rect 2692 4870 2722 4922
rect 2722 4870 2734 4922
rect 2734 4870 2748 4922
rect 2772 4870 2786 4922
rect 2786 4870 2798 4922
rect 2798 4870 2828 4922
rect 2852 4870 2862 4922
rect 2862 4870 2908 4922
rect 2612 4868 2668 4870
rect 2692 4868 2748 4870
rect 2772 4868 2828 4870
rect 2852 4868 2908 4870
rect 1214 4392 1270 4448
rect 2612 3834 2668 3836
rect 2692 3834 2748 3836
rect 2772 3834 2828 3836
rect 2852 3834 2908 3836
rect 2612 3782 2658 3834
rect 2658 3782 2668 3834
rect 2692 3782 2722 3834
rect 2722 3782 2734 3834
rect 2734 3782 2748 3834
rect 2772 3782 2786 3834
rect 2786 3782 2798 3834
rect 2798 3782 2828 3834
rect 2852 3782 2862 3834
rect 2862 3782 2908 3834
rect 2612 3780 2668 3782
rect 2692 3780 2748 3782
rect 2772 3780 2828 3782
rect 2852 3780 2908 3782
rect 1214 3304 1270 3360
rect 3348 5466 3404 5468
rect 3428 5466 3484 5468
rect 3508 5466 3564 5468
rect 3588 5466 3644 5468
rect 3348 5414 3394 5466
rect 3394 5414 3404 5466
rect 3428 5414 3458 5466
rect 3458 5414 3470 5466
rect 3470 5414 3484 5466
rect 3508 5414 3522 5466
rect 3522 5414 3534 5466
rect 3534 5414 3564 5466
rect 3588 5414 3598 5466
rect 3598 5414 3644 5466
rect 3348 5412 3404 5414
rect 3428 5412 3484 5414
rect 3508 5412 3564 5414
rect 3588 5412 3644 5414
rect 4820 6554 4876 6556
rect 4900 6554 4956 6556
rect 4980 6554 5036 6556
rect 5060 6554 5116 6556
rect 4820 6502 4866 6554
rect 4866 6502 4876 6554
rect 4900 6502 4930 6554
rect 4930 6502 4942 6554
rect 4942 6502 4956 6554
rect 4980 6502 4994 6554
rect 4994 6502 5006 6554
rect 5006 6502 5036 6554
rect 5060 6502 5070 6554
rect 5070 6502 5116 6554
rect 4820 6500 4876 6502
rect 4900 6500 4956 6502
rect 4980 6500 5036 6502
rect 5060 6500 5116 6502
rect 4084 6010 4140 6012
rect 4164 6010 4220 6012
rect 4244 6010 4300 6012
rect 4324 6010 4380 6012
rect 4084 5958 4130 6010
rect 4130 5958 4140 6010
rect 4164 5958 4194 6010
rect 4194 5958 4206 6010
rect 4206 5958 4220 6010
rect 4244 5958 4258 6010
rect 4258 5958 4270 6010
rect 4270 5958 4300 6010
rect 4324 5958 4334 6010
rect 4334 5958 4380 6010
rect 4084 5956 4140 5958
rect 4164 5956 4220 5958
rect 4244 5956 4300 5958
rect 4324 5956 4380 5958
rect 3348 4378 3404 4380
rect 3428 4378 3484 4380
rect 3508 4378 3564 4380
rect 3588 4378 3644 4380
rect 3348 4326 3394 4378
rect 3394 4326 3404 4378
rect 3428 4326 3458 4378
rect 3458 4326 3470 4378
rect 3470 4326 3484 4378
rect 3508 4326 3522 4378
rect 3522 4326 3534 4378
rect 3534 4326 3564 4378
rect 3588 4326 3598 4378
rect 3598 4326 3644 4378
rect 3348 4324 3404 4326
rect 3428 4324 3484 4326
rect 3508 4324 3564 4326
rect 3588 4324 3644 4326
rect 5556 7098 5612 7100
rect 5636 7098 5692 7100
rect 5716 7098 5772 7100
rect 5796 7098 5852 7100
rect 5556 7046 5602 7098
rect 5602 7046 5612 7098
rect 5636 7046 5666 7098
rect 5666 7046 5678 7098
rect 5678 7046 5692 7098
rect 5716 7046 5730 7098
rect 5730 7046 5742 7098
rect 5742 7046 5772 7098
rect 5796 7046 5806 7098
rect 5806 7046 5852 7098
rect 5556 7044 5612 7046
rect 5636 7044 5692 7046
rect 5716 7044 5772 7046
rect 5796 7044 5852 7046
rect 6292 6554 6348 6556
rect 6372 6554 6428 6556
rect 6452 6554 6508 6556
rect 6532 6554 6588 6556
rect 6292 6502 6338 6554
rect 6338 6502 6348 6554
rect 6372 6502 6402 6554
rect 6402 6502 6414 6554
rect 6414 6502 6428 6554
rect 6452 6502 6466 6554
rect 6466 6502 6478 6554
rect 6478 6502 6508 6554
rect 6532 6502 6542 6554
rect 6542 6502 6588 6554
rect 6292 6500 6348 6502
rect 6372 6500 6428 6502
rect 6452 6500 6508 6502
rect 6532 6500 6588 6502
rect 7028 7098 7084 7100
rect 7108 7098 7164 7100
rect 7188 7098 7244 7100
rect 7268 7098 7324 7100
rect 7028 7046 7074 7098
rect 7074 7046 7084 7098
rect 7108 7046 7138 7098
rect 7138 7046 7150 7098
rect 7150 7046 7164 7098
rect 7188 7046 7202 7098
rect 7202 7046 7214 7098
rect 7214 7046 7244 7098
rect 7268 7046 7278 7098
rect 7278 7046 7324 7098
rect 7028 7044 7084 7046
rect 7108 7044 7164 7046
rect 7188 7044 7244 7046
rect 7268 7044 7324 7046
rect 7764 7642 7820 7644
rect 7844 7642 7900 7644
rect 7924 7642 7980 7644
rect 8004 7642 8060 7644
rect 7764 7590 7810 7642
rect 7810 7590 7820 7642
rect 7844 7590 7874 7642
rect 7874 7590 7886 7642
rect 7886 7590 7900 7642
rect 7924 7590 7938 7642
rect 7938 7590 7950 7642
rect 7950 7590 7980 7642
rect 8004 7590 8014 7642
rect 8014 7590 8060 7642
rect 7764 7588 7820 7590
rect 7844 7588 7900 7590
rect 7924 7588 7980 7590
rect 8004 7588 8060 7590
rect 7764 6554 7820 6556
rect 7844 6554 7900 6556
rect 7924 6554 7980 6556
rect 8004 6554 8060 6556
rect 7764 6502 7810 6554
rect 7810 6502 7820 6554
rect 7844 6502 7874 6554
rect 7874 6502 7886 6554
rect 7886 6502 7900 6554
rect 7924 6502 7938 6554
rect 7938 6502 7950 6554
rect 7950 6502 7980 6554
rect 8004 6502 8014 6554
rect 8014 6502 8060 6554
rect 7764 6500 7820 6502
rect 7844 6500 7900 6502
rect 7924 6500 7980 6502
rect 8004 6500 8060 6502
rect 4084 4922 4140 4924
rect 4164 4922 4220 4924
rect 4244 4922 4300 4924
rect 4324 4922 4380 4924
rect 4084 4870 4130 4922
rect 4130 4870 4140 4922
rect 4164 4870 4194 4922
rect 4194 4870 4206 4922
rect 4206 4870 4220 4922
rect 4244 4870 4258 4922
rect 4258 4870 4270 4922
rect 4270 4870 4300 4922
rect 4324 4870 4334 4922
rect 4334 4870 4380 4922
rect 4084 4868 4140 4870
rect 4164 4868 4220 4870
rect 4244 4868 4300 4870
rect 4324 4868 4380 4870
rect 4084 3834 4140 3836
rect 4164 3834 4220 3836
rect 4244 3834 4300 3836
rect 4324 3834 4380 3836
rect 4084 3782 4130 3834
rect 4130 3782 4140 3834
rect 4164 3782 4194 3834
rect 4194 3782 4206 3834
rect 4206 3782 4220 3834
rect 4244 3782 4258 3834
rect 4258 3782 4270 3834
rect 4270 3782 4300 3834
rect 4324 3782 4334 3834
rect 4334 3782 4380 3834
rect 4084 3780 4140 3782
rect 4164 3780 4220 3782
rect 4244 3780 4300 3782
rect 4324 3780 4380 3782
rect 5556 6010 5612 6012
rect 5636 6010 5692 6012
rect 5716 6010 5772 6012
rect 5796 6010 5852 6012
rect 5556 5958 5602 6010
rect 5602 5958 5612 6010
rect 5636 5958 5666 6010
rect 5666 5958 5678 6010
rect 5678 5958 5692 6010
rect 5716 5958 5730 6010
rect 5730 5958 5742 6010
rect 5742 5958 5772 6010
rect 5796 5958 5806 6010
rect 5806 5958 5852 6010
rect 5556 5956 5612 5958
rect 5636 5956 5692 5958
rect 5716 5956 5772 5958
rect 5796 5956 5852 5958
rect 4820 5466 4876 5468
rect 4900 5466 4956 5468
rect 4980 5466 5036 5468
rect 5060 5466 5116 5468
rect 4820 5414 4866 5466
rect 4866 5414 4876 5466
rect 4900 5414 4930 5466
rect 4930 5414 4942 5466
rect 4942 5414 4956 5466
rect 4980 5414 4994 5466
rect 4994 5414 5006 5466
rect 5006 5414 5036 5466
rect 5060 5414 5070 5466
rect 5070 5414 5116 5466
rect 4820 5412 4876 5414
rect 4900 5412 4956 5414
rect 4980 5412 5036 5414
rect 5060 5412 5116 5414
rect 7028 6010 7084 6012
rect 7108 6010 7164 6012
rect 7188 6010 7244 6012
rect 7268 6010 7324 6012
rect 7028 5958 7074 6010
rect 7074 5958 7084 6010
rect 7108 5958 7138 6010
rect 7138 5958 7150 6010
rect 7150 5958 7164 6010
rect 7188 5958 7202 6010
rect 7202 5958 7214 6010
rect 7214 5958 7244 6010
rect 7268 5958 7278 6010
rect 7278 5958 7324 6010
rect 7028 5956 7084 5958
rect 7108 5956 7164 5958
rect 7188 5956 7244 5958
rect 7268 5956 7324 5958
rect 6292 5466 6348 5468
rect 6372 5466 6428 5468
rect 6452 5466 6508 5468
rect 6532 5466 6588 5468
rect 6292 5414 6338 5466
rect 6338 5414 6348 5466
rect 6372 5414 6402 5466
rect 6402 5414 6414 5466
rect 6414 5414 6428 5466
rect 6452 5414 6466 5466
rect 6466 5414 6478 5466
rect 6478 5414 6508 5466
rect 6532 5414 6542 5466
rect 6542 5414 6588 5466
rect 6292 5412 6348 5414
rect 6372 5412 6428 5414
rect 6452 5412 6508 5414
rect 6532 5412 6588 5414
rect 7764 5466 7820 5468
rect 7844 5466 7900 5468
rect 7924 5466 7980 5468
rect 8004 5466 8060 5468
rect 7764 5414 7810 5466
rect 7810 5414 7820 5466
rect 7844 5414 7874 5466
rect 7874 5414 7886 5466
rect 7886 5414 7900 5466
rect 7924 5414 7938 5466
rect 7938 5414 7950 5466
rect 7950 5414 7980 5466
rect 8004 5414 8014 5466
rect 8014 5414 8060 5466
rect 7764 5412 7820 5414
rect 7844 5412 7900 5414
rect 7924 5412 7980 5414
rect 8004 5412 8060 5414
rect 5556 4922 5612 4924
rect 5636 4922 5692 4924
rect 5716 4922 5772 4924
rect 5796 4922 5852 4924
rect 5556 4870 5602 4922
rect 5602 4870 5612 4922
rect 5636 4870 5666 4922
rect 5666 4870 5678 4922
rect 5678 4870 5692 4922
rect 5716 4870 5730 4922
rect 5730 4870 5742 4922
rect 5742 4870 5772 4922
rect 5796 4870 5806 4922
rect 5806 4870 5852 4922
rect 5556 4868 5612 4870
rect 5636 4868 5692 4870
rect 5716 4868 5772 4870
rect 5796 4868 5852 4870
rect 7028 4922 7084 4924
rect 7108 4922 7164 4924
rect 7188 4922 7244 4924
rect 7268 4922 7324 4924
rect 7028 4870 7074 4922
rect 7074 4870 7084 4922
rect 7108 4870 7138 4922
rect 7138 4870 7150 4922
rect 7150 4870 7164 4922
rect 7188 4870 7202 4922
rect 7202 4870 7214 4922
rect 7214 4870 7244 4922
rect 7268 4870 7278 4922
rect 7278 4870 7324 4922
rect 7028 4868 7084 4870
rect 7108 4868 7164 4870
rect 7188 4868 7244 4870
rect 7268 4868 7324 4870
rect 4820 4378 4876 4380
rect 4900 4378 4956 4380
rect 4980 4378 5036 4380
rect 5060 4378 5116 4380
rect 4820 4326 4866 4378
rect 4866 4326 4876 4378
rect 4900 4326 4930 4378
rect 4930 4326 4942 4378
rect 4942 4326 4956 4378
rect 4980 4326 4994 4378
rect 4994 4326 5006 4378
rect 5006 4326 5036 4378
rect 5060 4326 5070 4378
rect 5070 4326 5116 4378
rect 4820 4324 4876 4326
rect 4900 4324 4956 4326
rect 4980 4324 5036 4326
rect 5060 4324 5116 4326
rect 6292 4378 6348 4380
rect 6372 4378 6428 4380
rect 6452 4378 6508 4380
rect 6532 4378 6588 4380
rect 6292 4326 6338 4378
rect 6338 4326 6348 4378
rect 6372 4326 6402 4378
rect 6402 4326 6414 4378
rect 6414 4326 6428 4378
rect 6452 4326 6466 4378
rect 6466 4326 6478 4378
rect 6478 4326 6508 4378
rect 6532 4326 6542 4378
rect 6542 4326 6588 4378
rect 6292 4324 6348 4326
rect 6372 4324 6428 4326
rect 6452 4324 6508 4326
rect 6532 4324 6588 4326
rect 7764 4378 7820 4380
rect 7844 4378 7900 4380
rect 7924 4378 7980 4380
rect 8004 4378 8060 4380
rect 7764 4326 7810 4378
rect 7810 4326 7820 4378
rect 7844 4326 7874 4378
rect 7874 4326 7886 4378
rect 7886 4326 7900 4378
rect 7924 4326 7938 4378
rect 7938 4326 7950 4378
rect 7950 4326 7980 4378
rect 8004 4326 8014 4378
rect 8014 4326 8060 4378
rect 7764 4324 7820 4326
rect 7844 4324 7900 4326
rect 7924 4324 7980 4326
rect 8004 4324 8060 4326
rect 5556 3834 5612 3836
rect 5636 3834 5692 3836
rect 5716 3834 5772 3836
rect 5796 3834 5852 3836
rect 5556 3782 5602 3834
rect 5602 3782 5612 3834
rect 5636 3782 5666 3834
rect 5666 3782 5678 3834
rect 5678 3782 5692 3834
rect 5716 3782 5730 3834
rect 5730 3782 5742 3834
rect 5742 3782 5772 3834
rect 5796 3782 5806 3834
rect 5806 3782 5852 3834
rect 5556 3780 5612 3782
rect 5636 3780 5692 3782
rect 5716 3780 5772 3782
rect 5796 3780 5852 3782
rect 7028 3834 7084 3836
rect 7108 3834 7164 3836
rect 7188 3834 7244 3836
rect 7268 3834 7324 3836
rect 7028 3782 7074 3834
rect 7074 3782 7084 3834
rect 7108 3782 7138 3834
rect 7138 3782 7150 3834
rect 7150 3782 7164 3834
rect 7188 3782 7202 3834
rect 7202 3782 7214 3834
rect 7214 3782 7244 3834
rect 7268 3782 7278 3834
rect 7278 3782 7324 3834
rect 7028 3780 7084 3782
rect 7108 3780 7164 3782
rect 7188 3780 7244 3782
rect 7268 3780 7324 3782
rect 2612 2746 2668 2748
rect 2692 2746 2748 2748
rect 2772 2746 2828 2748
rect 2852 2746 2908 2748
rect 2612 2694 2658 2746
rect 2658 2694 2668 2746
rect 2692 2694 2722 2746
rect 2722 2694 2734 2746
rect 2734 2694 2748 2746
rect 2772 2694 2786 2746
rect 2786 2694 2798 2746
rect 2798 2694 2828 2746
rect 2852 2694 2862 2746
rect 2862 2694 2908 2746
rect 2612 2692 2668 2694
rect 2692 2692 2748 2694
rect 2772 2692 2828 2694
rect 2852 2692 2908 2694
rect 1214 2216 1270 2272
rect 3348 3290 3404 3292
rect 3428 3290 3484 3292
rect 3508 3290 3564 3292
rect 3588 3290 3644 3292
rect 3348 3238 3394 3290
rect 3394 3238 3404 3290
rect 3428 3238 3458 3290
rect 3458 3238 3470 3290
rect 3470 3238 3484 3290
rect 3508 3238 3522 3290
rect 3522 3238 3534 3290
rect 3534 3238 3564 3290
rect 3588 3238 3598 3290
rect 3598 3238 3644 3290
rect 3348 3236 3404 3238
rect 3428 3236 3484 3238
rect 3508 3236 3564 3238
rect 3588 3236 3644 3238
rect 4084 2746 4140 2748
rect 4164 2746 4220 2748
rect 4244 2746 4300 2748
rect 4324 2746 4380 2748
rect 4084 2694 4130 2746
rect 4130 2694 4140 2746
rect 4164 2694 4194 2746
rect 4194 2694 4206 2746
rect 4206 2694 4220 2746
rect 4244 2694 4258 2746
rect 4258 2694 4270 2746
rect 4270 2694 4300 2746
rect 4324 2694 4334 2746
rect 4334 2694 4380 2746
rect 4084 2692 4140 2694
rect 4164 2692 4220 2694
rect 4244 2692 4300 2694
rect 4324 2692 4380 2694
rect 4820 3290 4876 3292
rect 4900 3290 4956 3292
rect 4980 3290 5036 3292
rect 5060 3290 5116 3292
rect 4820 3238 4866 3290
rect 4866 3238 4876 3290
rect 4900 3238 4930 3290
rect 4930 3238 4942 3290
rect 4942 3238 4956 3290
rect 4980 3238 4994 3290
rect 4994 3238 5006 3290
rect 5006 3238 5036 3290
rect 5060 3238 5070 3290
rect 5070 3238 5116 3290
rect 4820 3236 4876 3238
rect 4900 3236 4956 3238
rect 4980 3236 5036 3238
rect 5060 3236 5116 3238
rect 6292 3290 6348 3292
rect 6372 3290 6428 3292
rect 6452 3290 6508 3292
rect 6532 3290 6588 3292
rect 6292 3238 6338 3290
rect 6338 3238 6348 3290
rect 6372 3238 6402 3290
rect 6402 3238 6414 3290
rect 6414 3238 6428 3290
rect 6452 3238 6466 3290
rect 6466 3238 6478 3290
rect 6478 3238 6508 3290
rect 6532 3238 6542 3290
rect 6542 3238 6588 3290
rect 6292 3236 6348 3238
rect 6372 3236 6428 3238
rect 6452 3236 6508 3238
rect 6532 3236 6588 3238
rect 5556 2746 5612 2748
rect 5636 2746 5692 2748
rect 5716 2746 5772 2748
rect 5796 2746 5852 2748
rect 5556 2694 5602 2746
rect 5602 2694 5612 2746
rect 5636 2694 5666 2746
rect 5666 2694 5678 2746
rect 5678 2694 5692 2746
rect 5716 2694 5730 2746
rect 5730 2694 5742 2746
rect 5742 2694 5772 2746
rect 5796 2694 5806 2746
rect 5806 2694 5852 2746
rect 5556 2692 5612 2694
rect 5636 2692 5692 2694
rect 5716 2692 5772 2694
rect 5796 2692 5852 2694
rect 7028 2746 7084 2748
rect 7108 2746 7164 2748
rect 7188 2746 7244 2748
rect 7268 2746 7324 2748
rect 7028 2694 7074 2746
rect 7074 2694 7084 2746
rect 7108 2694 7138 2746
rect 7138 2694 7150 2746
rect 7150 2694 7164 2746
rect 7188 2694 7202 2746
rect 7202 2694 7214 2746
rect 7214 2694 7244 2746
rect 7268 2694 7278 2746
rect 7278 2694 7324 2746
rect 7028 2692 7084 2694
rect 7108 2692 7164 2694
rect 7188 2692 7244 2694
rect 7268 2692 7324 2694
rect 7764 3290 7820 3292
rect 7844 3290 7900 3292
rect 7924 3290 7980 3292
rect 8004 3290 8060 3292
rect 7764 3238 7810 3290
rect 7810 3238 7820 3290
rect 7844 3238 7874 3290
rect 7874 3238 7886 3290
rect 7886 3238 7900 3290
rect 7924 3238 7938 3290
rect 7938 3238 7950 3290
rect 7950 3238 7980 3290
rect 8004 3238 8014 3290
rect 8014 3238 8060 3290
rect 7764 3236 7820 3238
rect 7844 3236 7900 3238
rect 7924 3236 7980 3238
rect 8004 3236 8060 3238
rect 3348 2202 3404 2204
rect 3428 2202 3484 2204
rect 3508 2202 3564 2204
rect 3588 2202 3644 2204
rect 3348 2150 3394 2202
rect 3394 2150 3404 2202
rect 3428 2150 3458 2202
rect 3458 2150 3470 2202
rect 3470 2150 3484 2202
rect 3508 2150 3522 2202
rect 3522 2150 3534 2202
rect 3534 2150 3564 2202
rect 3588 2150 3598 2202
rect 3598 2150 3644 2202
rect 3348 2148 3404 2150
rect 3428 2148 3484 2150
rect 3508 2148 3564 2150
rect 3588 2148 3644 2150
rect 4820 2202 4876 2204
rect 4900 2202 4956 2204
rect 4980 2202 5036 2204
rect 5060 2202 5116 2204
rect 4820 2150 4866 2202
rect 4866 2150 4876 2202
rect 4900 2150 4930 2202
rect 4930 2150 4942 2202
rect 4942 2150 4956 2202
rect 4980 2150 4994 2202
rect 4994 2150 5006 2202
rect 5006 2150 5036 2202
rect 5060 2150 5070 2202
rect 5070 2150 5116 2202
rect 4820 2148 4876 2150
rect 4900 2148 4956 2150
rect 4980 2148 5036 2150
rect 5060 2148 5116 2150
rect 6292 2202 6348 2204
rect 6372 2202 6428 2204
rect 6452 2202 6508 2204
rect 6532 2202 6588 2204
rect 6292 2150 6338 2202
rect 6338 2150 6348 2202
rect 6372 2150 6402 2202
rect 6402 2150 6414 2202
rect 6414 2150 6428 2202
rect 6452 2150 6466 2202
rect 6466 2150 6478 2202
rect 6478 2150 6508 2202
rect 6532 2150 6542 2202
rect 6542 2150 6588 2202
rect 6292 2148 6348 2150
rect 6372 2148 6428 2150
rect 6452 2148 6508 2150
rect 6532 2148 6588 2150
rect 7764 2202 7820 2204
rect 7844 2202 7900 2204
rect 7924 2202 7980 2204
rect 8004 2202 8060 2204
rect 7764 2150 7810 2202
rect 7810 2150 7820 2202
rect 7844 2150 7874 2202
rect 7874 2150 7886 2202
rect 7886 2150 7900 2202
rect 7924 2150 7938 2202
rect 7938 2150 7950 2202
rect 7950 2150 7980 2202
rect 8004 2150 8014 2202
rect 8014 2150 8060 2202
rect 7764 2148 7820 2150
rect 7844 2148 7900 2150
rect 7924 2148 7980 2150
rect 8004 2148 8060 2150
rect 3054 1128 3110 1184
<< metal3 >>
rect 0 8802 400 8832
rect 2957 8802 3023 8805
rect 0 8800 3023 8802
rect 0 8744 2962 8800
rect 3018 8744 3023 8800
rect 0 8742 3023 8744
rect 0 8712 400 8742
rect 2957 8739 3023 8742
rect 0 7714 400 7744
rect 841 7714 907 7717
rect 0 7712 907 7714
rect 0 7656 846 7712
rect 902 7656 907 7712
rect 0 7654 907 7656
rect 0 7624 400 7654
rect 841 7651 907 7654
rect 3338 7648 3654 7649
rect 3338 7584 3344 7648
rect 3408 7584 3424 7648
rect 3488 7584 3504 7648
rect 3568 7584 3584 7648
rect 3648 7584 3654 7648
rect 3338 7583 3654 7584
rect 4810 7648 5126 7649
rect 4810 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5126 7648
rect 4810 7583 5126 7584
rect 6282 7648 6598 7649
rect 6282 7584 6288 7648
rect 6352 7584 6368 7648
rect 6432 7584 6448 7648
rect 6512 7584 6528 7648
rect 6592 7584 6598 7648
rect 6282 7583 6598 7584
rect 7754 7648 8070 7649
rect 7754 7584 7760 7648
rect 7824 7584 7840 7648
rect 7904 7584 7920 7648
rect 7984 7584 8000 7648
rect 8064 7584 8070 7648
rect 7754 7583 8070 7584
rect 2602 7104 2918 7105
rect 2602 7040 2608 7104
rect 2672 7040 2688 7104
rect 2752 7040 2768 7104
rect 2832 7040 2848 7104
rect 2912 7040 2918 7104
rect 2602 7039 2918 7040
rect 4074 7104 4390 7105
rect 4074 7040 4080 7104
rect 4144 7040 4160 7104
rect 4224 7040 4240 7104
rect 4304 7040 4320 7104
rect 4384 7040 4390 7104
rect 4074 7039 4390 7040
rect 5546 7104 5862 7105
rect 5546 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5862 7104
rect 5546 7039 5862 7040
rect 7018 7104 7334 7105
rect 7018 7040 7024 7104
rect 7088 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7334 7104
rect 7018 7039 7334 7040
rect 0 6626 400 6656
rect 1301 6626 1367 6629
rect 0 6624 1367 6626
rect 0 6568 1306 6624
rect 1362 6568 1367 6624
rect 0 6566 1367 6568
rect 0 6536 400 6566
rect 1301 6563 1367 6566
rect 3338 6560 3654 6561
rect 3338 6496 3344 6560
rect 3408 6496 3424 6560
rect 3488 6496 3504 6560
rect 3568 6496 3584 6560
rect 3648 6496 3654 6560
rect 3338 6495 3654 6496
rect 4810 6560 5126 6561
rect 4810 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5126 6560
rect 4810 6495 5126 6496
rect 6282 6560 6598 6561
rect 6282 6496 6288 6560
rect 6352 6496 6368 6560
rect 6432 6496 6448 6560
rect 6512 6496 6528 6560
rect 6592 6496 6598 6560
rect 6282 6495 6598 6496
rect 7754 6560 8070 6561
rect 7754 6496 7760 6560
rect 7824 6496 7840 6560
rect 7904 6496 7920 6560
rect 7984 6496 8000 6560
rect 8064 6496 8070 6560
rect 7754 6495 8070 6496
rect 2602 6016 2918 6017
rect 2602 5952 2608 6016
rect 2672 5952 2688 6016
rect 2752 5952 2768 6016
rect 2832 5952 2848 6016
rect 2912 5952 2918 6016
rect 2602 5951 2918 5952
rect 4074 6016 4390 6017
rect 4074 5952 4080 6016
rect 4144 5952 4160 6016
rect 4224 5952 4240 6016
rect 4304 5952 4320 6016
rect 4384 5952 4390 6016
rect 4074 5951 4390 5952
rect 5546 6016 5862 6017
rect 5546 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5862 6016
rect 5546 5951 5862 5952
rect 7018 6016 7334 6017
rect 7018 5952 7024 6016
rect 7088 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7334 6016
rect 7018 5951 7334 5952
rect 0 5538 400 5568
rect 2405 5538 2471 5541
rect 0 5536 2471 5538
rect 0 5480 2410 5536
rect 2466 5480 2471 5536
rect 0 5478 2471 5480
rect 0 5448 400 5478
rect 2405 5475 2471 5478
rect 3338 5472 3654 5473
rect 3338 5408 3344 5472
rect 3408 5408 3424 5472
rect 3488 5408 3504 5472
rect 3568 5408 3584 5472
rect 3648 5408 3654 5472
rect 3338 5407 3654 5408
rect 4810 5472 5126 5473
rect 4810 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5126 5472
rect 4810 5407 5126 5408
rect 6282 5472 6598 5473
rect 6282 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6598 5472
rect 6282 5407 6598 5408
rect 7754 5472 8070 5473
rect 7754 5408 7760 5472
rect 7824 5408 7840 5472
rect 7904 5408 7920 5472
rect 7984 5408 8000 5472
rect 8064 5408 8070 5472
rect 7754 5407 8070 5408
rect 2602 4928 2918 4929
rect 2602 4864 2608 4928
rect 2672 4864 2688 4928
rect 2752 4864 2768 4928
rect 2832 4864 2848 4928
rect 2912 4864 2918 4928
rect 2602 4863 2918 4864
rect 4074 4928 4390 4929
rect 4074 4864 4080 4928
rect 4144 4864 4160 4928
rect 4224 4864 4240 4928
rect 4304 4864 4320 4928
rect 4384 4864 4390 4928
rect 4074 4863 4390 4864
rect 5546 4928 5862 4929
rect 5546 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5862 4928
rect 5546 4863 5862 4864
rect 7018 4928 7334 4929
rect 7018 4864 7024 4928
rect 7088 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7334 4928
rect 7018 4863 7334 4864
rect 0 4450 400 4480
rect 1209 4450 1275 4453
rect 0 4448 1275 4450
rect 0 4392 1214 4448
rect 1270 4392 1275 4448
rect 0 4390 1275 4392
rect 0 4360 400 4390
rect 1209 4387 1275 4390
rect 3338 4384 3654 4385
rect 3338 4320 3344 4384
rect 3408 4320 3424 4384
rect 3488 4320 3504 4384
rect 3568 4320 3584 4384
rect 3648 4320 3654 4384
rect 3338 4319 3654 4320
rect 4810 4384 5126 4385
rect 4810 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5126 4384
rect 4810 4319 5126 4320
rect 6282 4384 6598 4385
rect 6282 4320 6288 4384
rect 6352 4320 6368 4384
rect 6432 4320 6448 4384
rect 6512 4320 6528 4384
rect 6592 4320 6598 4384
rect 6282 4319 6598 4320
rect 7754 4384 8070 4385
rect 7754 4320 7760 4384
rect 7824 4320 7840 4384
rect 7904 4320 7920 4384
rect 7984 4320 8000 4384
rect 8064 4320 8070 4384
rect 7754 4319 8070 4320
rect 2602 3840 2918 3841
rect 2602 3776 2608 3840
rect 2672 3776 2688 3840
rect 2752 3776 2768 3840
rect 2832 3776 2848 3840
rect 2912 3776 2918 3840
rect 2602 3775 2918 3776
rect 4074 3840 4390 3841
rect 4074 3776 4080 3840
rect 4144 3776 4160 3840
rect 4224 3776 4240 3840
rect 4304 3776 4320 3840
rect 4384 3776 4390 3840
rect 4074 3775 4390 3776
rect 5546 3840 5862 3841
rect 5546 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5862 3840
rect 5546 3775 5862 3776
rect 7018 3840 7334 3841
rect 7018 3776 7024 3840
rect 7088 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7334 3840
rect 7018 3775 7334 3776
rect 0 3362 400 3392
rect 1209 3362 1275 3365
rect 0 3360 1275 3362
rect 0 3304 1214 3360
rect 1270 3304 1275 3360
rect 0 3302 1275 3304
rect 0 3272 400 3302
rect 1209 3299 1275 3302
rect 3338 3296 3654 3297
rect 3338 3232 3344 3296
rect 3408 3232 3424 3296
rect 3488 3232 3504 3296
rect 3568 3232 3584 3296
rect 3648 3232 3654 3296
rect 3338 3231 3654 3232
rect 4810 3296 5126 3297
rect 4810 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5126 3296
rect 4810 3231 5126 3232
rect 6282 3296 6598 3297
rect 6282 3232 6288 3296
rect 6352 3232 6368 3296
rect 6432 3232 6448 3296
rect 6512 3232 6528 3296
rect 6592 3232 6598 3296
rect 6282 3231 6598 3232
rect 7754 3296 8070 3297
rect 7754 3232 7760 3296
rect 7824 3232 7840 3296
rect 7904 3232 7920 3296
rect 7984 3232 8000 3296
rect 8064 3232 8070 3296
rect 7754 3231 8070 3232
rect 2602 2752 2918 2753
rect 2602 2688 2608 2752
rect 2672 2688 2688 2752
rect 2752 2688 2768 2752
rect 2832 2688 2848 2752
rect 2912 2688 2918 2752
rect 2602 2687 2918 2688
rect 4074 2752 4390 2753
rect 4074 2688 4080 2752
rect 4144 2688 4160 2752
rect 4224 2688 4240 2752
rect 4304 2688 4320 2752
rect 4384 2688 4390 2752
rect 4074 2687 4390 2688
rect 5546 2752 5862 2753
rect 5546 2688 5552 2752
rect 5616 2688 5632 2752
rect 5696 2688 5712 2752
rect 5776 2688 5792 2752
rect 5856 2688 5862 2752
rect 5546 2687 5862 2688
rect 7018 2752 7334 2753
rect 7018 2688 7024 2752
rect 7088 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7334 2752
rect 7018 2687 7334 2688
rect 0 2274 400 2304
rect 1209 2274 1275 2277
rect 0 2272 1275 2274
rect 0 2216 1214 2272
rect 1270 2216 1275 2272
rect 0 2214 1275 2216
rect 0 2184 400 2214
rect 1209 2211 1275 2214
rect 3338 2208 3654 2209
rect 3338 2144 3344 2208
rect 3408 2144 3424 2208
rect 3488 2144 3504 2208
rect 3568 2144 3584 2208
rect 3648 2144 3654 2208
rect 3338 2143 3654 2144
rect 4810 2208 5126 2209
rect 4810 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5126 2208
rect 4810 2143 5126 2144
rect 6282 2208 6598 2209
rect 6282 2144 6288 2208
rect 6352 2144 6368 2208
rect 6432 2144 6448 2208
rect 6512 2144 6528 2208
rect 6592 2144 6598 2208
rect 6282 2143 6598 2144
rect 7754 2208 8070 2209
rect 7754 2144 7760 2208
rect 7824 2144 7840 2208
rect 7904 2144 7920 2208
rect 7984 2144 8000 2208
rect 8064 2144 8070 2208
rect 7754 2143 8070 2144
rect 0 1186 400 1216
rect 3049 1186 3115 1189
rect 0 1184 3115 1186
rect 0 1128 3054 1184
rect 3110 1128 3115 1184
rect 0 1126 3115 1128
rect 0 1096 400 1126
rect 3049 1123 3115 1126
<< via3 >>
rect 3344 7644 3408 7648
rect 3344 7588 3348 7644
rect 3348 7588 3404 7644
rect 3404 7588 3408 7644
rect 3344 7584 3408 7588
rect 3424 7644 3488 7648
rect 3424 7588 3428 7644
rect 3428 7588 3484 7644
rect 3484 7588 3488 7644
rect 3424 7584 3488 7588
rect 3504 7644 3568 7648
rect 3504 7588 3508 7644
rect 3508 7588 3564 7644
rect 3564 7588 3568 7644
rect 3504 7584 3568 7588
rect 3584 7644 3648 7648
rect 3584 7588 3588 7644
rect 3588 7588 3644 7644
rect 3644 7588 3648 7644
rect 3584 7584 3648 7588
rect 4816 7644 4880 7648
rect 4816 7588 4820 7644
rect 4820 7588 4876 7644
rect 4876 7588 4880 7644
rect 4816 7584 4880 7588
rect 4896 7644 4960 7648
rect 4896 7588 4900 7644
rect 4900 7588 4956 7644
rect 4956 7588 4960 7644
rect 4896 7584 4960 7588
rect 4976 7644 5040 7648
rect 4976 7588 4980 7644
rect 4980 7588 5036 7644
rect 5036 7588 5040 7644
rect 4976 7584 5040 7588
rect 5056 7644 5120 7648
rect 5056 7588 5060 7644
rect 5060 7588 5116 7644
rect 5116 7588 5120 7644
rect 5056 7584 5120 7588
rect 6288 7644 6352 7648
rect 6288 7588 6292 7644
rect 6292 7588 6348 7644
rect 6348 7588 6352 7644
rect 6288 7584 6352 7588
rect 6368 7644 6432 7648
rect 6368 7588 6372 7644
rect 6372 7588 6428 7644
rect 6428 7588 6432 7644
rect 6368 7584 6432 7588
rect 6448 7644 6512 7648
rect 6448 7588 6452 7644
rect 6452 7588 6508 7644
rect 6508 7588 6512 7644
rect 6448 7584 6512 7588
rect 6528 7644 6592 7648
rect 6528 7588 6532 7644
rect 6532 7588 6588 7644
rect 6588 7588 6592 7644
rect 6528 7584 6592 7588
rect 7760 7644 7824 7648
rect 7760 7588 7764 7644
rect 7764 7588 7820 7644
rect 7820 7588 7824 7644
rect 7760 7584 7824 7588
rect 7840 7644 7904 7648
rect 7840 7588 7844 7644
rect 7844 7588 7900 7644
rect 7900 7588 7904 7644
rect 7840 7584 7904 7588
rect 7920 7644 7984 7648
rect 7920 7588 7924 7644
rect 7924 7588 7980 7644
rect 7980 7588 7984 7644
rect 7920 7584 7984 7588
rect 8000 7644 8064 7648
rect 8000 7588 8004 7644
rect 8004 7588 8060 7644
rect 8060 7588 8064 7644
rect 8000 7584 8064 7588
rect 2608 7100 2672 7104
rect 2608 7044 2612 7100
rect 2612 7044 2668 7100
rect 2668 7044 2672 7100
rect 2608 7040 2672 7044
rect 2688 7100 2752 7104
rect 2688 7044 2692 7100
rect 2692 7044 2748 7100
rect 2748 7044 2752 7100
rect 2688 7040 2752 7044
rect 2768 7100 2832 7104
rect 2768 7044 2772 7100
rect 2772 7044 2828 7100
rect 2828 7044 2832 7100
rect 2768 7040 2832 7044
rect 2848 7100 2912 7104
rect 2848 7044 2852 7100
rect 2852 7044 2908 7100
rect 2908 7044 2912 7100
rect 2848 7040 2912 7044
rect 4080 7100 4144 7104
rect 4080 7044 4084 7100
rect 4084 7044 4140 7100
rect 4140 7044 4144 7100
rect 4080 7040 4144 7044
rect 4160 7100 4224 7104
rect 4160 7044 4164 7100
rect 4164 7044 4220 7100
rect 4220 7044 4224 7100
rect 4160 7040 4224 7044
rect 4240 7100 4304 7104
rect 4240 7044 4244 7100
rect 4244 7044 4300 7100
rect 4300 7044 4304 7100
rect 4240 7040 4304 7044
rect 4320 7100 4384 7104
rect 4320 7044 4324 7100
rect 4324 7044 4380 7100
rect 4380 7044 4384 7100
rect 4320 7040 4384 7044
rect 5552 7100 5616 7104
rect 5552 7044 5556 7100
rect 5556 7044 5612 7100
rect 5612 7044 5616 7100
rect 5552 7040 5616 7044
rect 5632 7100 5696 7104
rect 5632 7044 5636 7100
rect 5636 7044 5692 7100
rect 5692 7044 5696 7100
rect 5632 7040 5696 7044
rect 5712 7100 5776 7104
rect 5712 7044 5716 7100
rect 5716 7044 5772 7100
rect 5772 7044 5776 7100
rect 5712 7040 5776 7044
rect 5792 7100 5856 7104
rect 5792 7044 5796 7100
rect 5796 7044 5852 7100
rect 5852 7044 5856 7100
rect 5792 7040 5856 7044
rect 7024 7100 7088 7104
rect 7024 7044 7028 7100
rect 7028 7044 7084 7100
rect 7084 7044 7088 7100
rect 7024 7040 7088 7044
rect 7104 7100 7168 7104
rect 7104 7044 7108 7100
rect 7108 7044 7164 7100
rect 7164 7044 7168 7100
rect 7104 7040 7168 7044
rect 7184 7100 7248 7104
rect 7184 7044 7188 7100
rect 7188 7044 7244 7100
rect 7244 7044 7248 7100
rect 7184 7040 7248 7044
rect 7264 7100 7328 7104
rect 7264 7044 7268 7100
rect 7268 7044 7324 7100
rect 7324 7044 7328 7100
rect 7264 7040 7328 7044
rect 3344 6556 3408 6560
rect 3344 6500 3348 6556
rect 3348 6500 3404 6556
rect 3404 6500 3408 6556
rect 3344 6496 3408 6500
rect 3424 6556 3488 6560
rect 3424 6500 3428 6556
rect 3428 6500 3484 6556
rect 3484 6500 3488 6556
rect 3424 6496 3488 6500
rect 3504 6556 3568 6560
rect 3504 6500 3508 6556
rect 3508 6500 3564 6556
rect 3564 6500 3568 6556
rect 3504 6496 3568 6500
rect 3584 6556 3648 6560
rect 3584 6500 3588 6556
rect 3588 6500 3644 6556
rect 3644 6500 3648 6556
rect 3584 6496 3648 6500
rect 4816 6556 4880 6560
rect 4816 6500 4820 6556
rect 4820 6500 4876 6556
rect 4876 6500 4880 6556
rect 4816 6496 4880 6500
rect 4896 6556 4960 6560
rect 4896 6500 4900 6556
rect 4900 6500 4956 6556
rect 4956 6500 4960 6556
rect 4896 6496 4960 6500
rect 4976 6556 5040 6560
rect 4976 6500 4980 6556
rect 4980 6500 5036 6556
rect 5036 6500 5040 6556
rect 4976 6496 5040 6500
rect 5056 6556 5120 6560
rect 5056 6500 5060 6556
rect 5060 6500 5116 6556
rect 5116 6500 5120 6556
rect 5056 6496 5120 6500
rect 6288 6556 6352 6560
rect 6288 6500 6292 6556
rect 6292 6500 6348 6556
rect 6348 6500 6352 6556
rect 6288 6496 6352 6500
rect 6368 6556 6432 6560
rect 6368 6500 6372 6556
rect 6372 6500 6428 6556
rect 6428 6500 6432 6556
rect 6368 6496 6432 6500
rect 6448 6556 6512 6560
rect 6448 6500 6452 6556
rect 6452 6500 6508 6556
rect 6508 6500 6512 6556
rect 6448 6496 6512 6500
rect 6528 6556 6592 6560
rect 6528 6500 6532 6556
rect 6532 6500 6588 6556
rect 6588 6500 6592 6556
rect 6528 6496 6592 6500
rect 7760 6556 7824 6560
rect 7760 6500 7764 6556
rect 7764 6500 7820 6556
rect 7820 6500 7824 6556
rect 7760 6496 7824 6500
rect 7840 6556 7904 6560
rect 7840 6500 7844 6556
rect 7844 6500 7900 6556
rect 7900 6500 7904 6556
rect 7840 6496 7904 6500
rect 7920 6556 7984 6560
rect 7920 6500 7924 6556
rect 7924 6500 7980 6556
rect 7980 6500 7984 6556
rect 7920 6496 7984 6500
rect 8000 6556 8064 6560
rect 8000 6500 8004 6556
rect 8004 6500 8060 6556
rect 8060 6500 8064 6556
rect 8000 6496 8064 6500
rect 2608 6012 2672 6016
rect 2608 5956 2612 6012
rect 2612 5956 2668 6012
rect 2668 5956 2672 6012
rect 2608 5952 2672 5956
rect 2688 6012 2752 6016
rect 2688 5956 2692 6012
rect 2692 5956 2748 6012
rect 2748 5956 2752 6012
rect 2688 5952 2752 5956
rect 2768 6012 2832 6016
rect 2768 5956 2772 6012
rect 2772 5956 2828 6012
rect 2828 5956 2832 6012
rect 2768 5952 2832 5956
rect 2848 6012 2912 6016
rect 2848 5956 2852 6012
rect 2852 5956 2908 6012
rect 2908 5956 2912 6012
rect 2848 5952 2912 5956
rect 4080 6012 4144 6016
rect 4080 5956 4084 6012
rect 4084 5956 4140 6012
rect 4140 5956 4144 6012
rect 4080 5952 4144 5956
rect 4160 6012 4224 6016
rect 4160 5956 4164 6012
rect 4164 5956 4220 6012
rect 4220 5956 4224 6012
rect 4160 5952 4224 5956
rect 4240 6012 4304 6016
rect 4240 5956 4244 6012
rect 4244 5956 4300 6012
rect 4300 5956 4304 6012
rect 4240 5952 4304 5956
rect 4320 6012 4384 6016
rect 4320 5956 4324 6012
rect 4324 5956 4380 6012
rect 4380 5956 4384 6012
rect 4320 5952 4384 5956
rect 5552 6012 5616 6016
rect 5552 5956 5556 6012
rect 5556 5956 5612 6012
rect 5612 5956 5616 6012
rect 5552 5952 5616 5956
rect 5632 6012 5696 6016
rect 5632 5956 5636 6012
rect 5636 5956 5692 6012
rect 5692 5956 5696 6012
rect 5632 5952 5696 5956
rect 5712 6012 5776 6016
rect 5712 5956 5716 6012
rect 5716 5956 5772 6012
rect 5772 5956 5776 6012
rect 5712 5952 5776 5956
rect 5792 6012 5856 6016
rect 5792 5956 5796 6012
rect 5796 5956 5852 6012
rect 5852 5956 5856 6012
rect 5792 5952 5856 5956
rect 7024 6012 7088 6016
rect 7024 5956 7028 6012
rect 7028 5956 7084 6012
rect 7084 5956 7088 6012
rect 7024 5952 7088 5956
rect 7104 6012 7168 6016
rect 7104 5956 7108 6012
rect 7108 5956 7164 6012
rect 7164 5956 7168 6012
rect 7104 5952 7168 5956
rect 7184 6012 7248 6016
rect 7184 5956 7188 6012
rect 7188 5956 7244 6012
rect 7244 5956 7248 6012
rect 7184 5952 7248 5956
rect 7264 6012 7328 6016
rect 7264 5956 7268 6012
rect 7268 5956 7324 6012
rect 7324 5956 7328 6012
rect 7264 5952 7328 5956
rect 3344 5468 3408 5472
rect 3344 5412 3348 5468
rect 3348 5412 3404 5468
rect 3404 5412 3408 5468
rect 3344 5408 3408 5412
rect 3424 5468 3488 5472
rect 3424 5412 3428 5468
rect 3428 5412 3484 5468
rect 3484 5412 3488 5468
rect 3424 5408 3488 5412
rect 3504 5468 3568 5472
rect 3504 5412 3508 5468
rect 3508 5412 3564 5468
rect 3564 5412 3568 5468
rect 3504 5408 3568 5412
rect 3584 5468 3648 5472
rect 3584 5412 3588 5468
rect 3588 5412 3644 5468
rect 3644 5412 3648 5468
rect 3584 5408 3648 5412
rect 4816 5468 4880 5472
rect 4816 5412 4820 5468
rect 4820 5412 4876 5468
rect 4876 5412 4880 5468
rect 4816 5408 4880 5412
rect 4896 5468 4960 5472
rect 4896 5412 4900 5468
rect 4900 5412 4956 5468
rect 4956 5412 4960 5468
rect 4896 5408 4960 5412
rect 4976 5468 5040 5472
rect 4976 5412 4980 5468
rect 4980 5412 5036 5468
rect 5036 5412 5040 5468
rect 4976 5408 5040 5412
rect 5056 5468 5120 5472
rect 5056 5412 5060 5468
rect 5060 5412 5116 5468
rect 5116 5412 5120 5468
rect 5056 5408 5120 5412
rect 6288 5468 6352 5472
rect 6288 5412 6292 5468
rect 6292 5412 6348 5468
rect 6348 5412 6352 5468
rect 6288 5408 6352 5412
rect 6368 5468 6432 5472
rect 6368 5412 6372 5468
rect 6372 5412 6428 5468
rect 6428 5412 6432 5468
rect 6368 5408 6432 5412
rect 6448 5468 6512 5472
rect 6448 5412 6452 5468
rect 6452 5412 6508 5468
rect 6508 5412 6512 5468
rect 6448 5408 6512 5412
rect 6528 5468 6592 5472
rect 6528 5412 6532 5468
rect 6532 5412 6588 5468
rect 6588 5412 6592 5468
rect 6528 5408 6592 5412
rect 7760 5468 7824 5472
rect 7760 5412 7764 5468
rect 7764 5412 7820 5468
rect 7820 5412 7824 5468
rect 7760 5408 7824 5412
rect 7840 5468 7904 5472
rect 7840 5412 7844 5468
rect 7844 5412 7900 5468
rect 7900 5412 7904 5468
rect 7840 5408 7904 5412
rect 7920 5468 7984 5472
rect 7920 5412 7924 5468
rect 7924 5412 7980 5468
rect 7980 5412 7984 5468
rect 7920 5408 7984 5412
rect 8000 5468 8064 5472
rect 8000 5412 8004 5468
rect 8004 5412 8060 5468
rect 8060 5412 8064 5468
rect 8000 5408 8064 5412
rect 2608 4924 2672 4928
rect 2608 4868 2612 4924
rect 2612 4868 2668 4924
rect 2668 4868 2672 4924
rect 2608 4864 2672 4868
rect 2688 4924 2752 4928
rect 2688 4868 2692 4924
rect 2692 4868 2748 4924
rect 2748 4868 2752 4924
rect 2688 4864 2752 4868
rect 2768 4924 2832 4928
rect 2768 4868 2772 4924
rect 2772 4868 2828 4924
rect 2828 4868 2832 4924
rect 2768 4864 2832 4868
rect 2848 4924 2912 4928
rect 2848 4868 2852 4924
rect 2852 4868 2908 4924
rect 2908 4868 2912 4924
rect 2848 4864 2912 4868
rect 4080 4924 4144 4928
rect 4080 4868 4084 4924
rect 4084 4868 4140 4924
rect 4140 4868 4144 4924
rect 4080 4864 4144 4868
rect 4160 4924 4224 4928
rect 4160 4868 4164 4924
rect 4164 4868 4220 4924
rect 4220 4868 4224 4924
rect 4160 4864 4224 4868
rect 4240 4924 4304 4928
rect 4240 4868 4244 4924
rect 4244 4868 4300 4924
rect 4300 4868 4304 4924
rect 4240 4864 4304 4868
rect 4320 4924 4384 4928
rect 4320 4868 4324 4924
rect 4324 4868 4380 4924
rect 4380 4868 4384 4924
rect 4320 4864 4384 4868
rect 5552 4924 5616 4928
rect 5552 4868 5556 4924
rect 5556 4868 5612 4924
rect 5612 4868 5616 4924
rect 5552 4864 5616 4868
rect 5632 4924 5696 4928
rect 5632 4868 5636 4924
rect 5636 4868 5692 4924
rect 5692 4868 5696 4924
rect 5632 4864 5696 4868
rect 5712 4924 5776 4928
rect 5712 4868 5716 4924
rect 5716 4868 5772 4924
rect 5772 4868 5776 4924
rect 5712 4864 5776 4868
rect 5792 4924 5856 4928
rect 5792 4868 5796 4924
rect 5796 4868 5852 4924
rect 5852 4868 5856 4924
rect 5792 4864 5856 4868
rect 7024 4924 7088 4928
rect 7024 4868 7028 4924
rect 7028 4868 7084 4924
rect 7084 4868 7088 4924
rect 7024 4864 7088 4868
rect 7104 4924 7168 4928
rect 7104 4868 7108 4924
rect 7108 4868 7164 4924
rect 7164 4868 7168 4924
rect 7104 4864 7168 4868
rect 7184 4924 7248 4928
rect 7184 4868 7188 4924
rect 7188 4868 7244 4924
rect 7244 4868 7248 4924
rect 7184 4864 7248 4868
rect 7264 4924 7328 4928
rect 7264 4868 7268 4924
rect 7268 4868 7324 4924
rect 7324 4868 7328 4924
rect 7264 4864 7328 4868
rect 3344 4380 3408 4384
rect 3344 4324 3348 4380
rect 3348 4324 3404 4380
rect 3404 4324 3408 4380
rect 3344 4320 3408 4324
rect 3424 4380 3488 4384
rect 3424 4324 3428 4380
rect 3428 4324 3484 4380
rect 3484 4324 3488 4380
rect 3424 4320 3488 4324
rect 3504 4380 3568 4384
rect 3504 4324 3508 4380
rect 3508 4324 3564 4380
rect 3564 4324 3568 4380
rect 3504 4320 3568 4324
rect 3584 4380 3648 4384
rect 3584 4324 3588 4380
rect 3588 4324 3644 4380
rect 3644 4324 3648 4380
rect 3584 4320 3648 4324
rect 4816 4380 4880 4384
rect 4816 4324 4820 4380
rect 4820 4324 4876 4380
rect 4876 4324 4880 4380
rect 4816 4320 4880 4324
rect 4896 4380 4960 4384
rect 4896 4324 4900 4380
rect 4900 4324 4956 4380
rect 4956 4324 4960 4380
rect 4896 4320 4960 4324
rect 4976 4380 5040 4384
rect 4976 4324 4980 4380
rect 4980 4324 5036 4380
rect 5036 4324 5040 4380
rect 4976 4320 5040 4324
rect 5056 4380 5120 4384
rect 5056 4324 5060 4380
rect 5060 4324 5116 4380
rect 5116 4324 5120 4380
rect 5056 4320 5120 4324
rect 6288 4380 6352 4384
rect 6288 4324 6292 4380
rect 6292 4324 6348 4380
rect 6348 4324 6352 4380
rect 6288 4320 6352 4324
rect 6368 4380 6432 4384
rect 6368 4324 6372 4380
rect 6372 4324 6428 4380
rect 6428 4324 6432 4380
rect 6368 4320 6432 4324
rect 6448 4380 6512 4384
rect 6448 4324 6452 4380
rect 6452 4324 6508 4380
rect 6508 4324 6512 4380
rect 6448 4320 6512 4324
rect 6528 4380 6592 4384
rect 6528 4324 6532 4380
rect 6532 4324 6588 4380
rect 6588 4324 6592 4380
rect 6528 4320 6592 4324
rect 7760 4380 7824 4384
rect 7760 4324 7764 4380
rect 7764 4324 7820 4380
rect 7820 4324 7824 4380
rect 7760 4320 7824 4324
rect 7840 4380 7904 4384
rect 7840 4324 7844 4380
rect 7844 4324 7900 4380
rect 7900 4324 7904 4380
rect 7840 4320 7904 4324
rect 7920 4380 7984 4384
rect 7920 4324 7924 4380
rect 7924 4324 7980 4380
rect 7980 4324 7984 4380
rect 7920 4320 7984 4324
rect 8000 4380 8064 4384
rect 8000 4324 8004 4380
rect 8004 4324 8060 4380
rect 8060 4324 8064 4380
rect 8000 4320 8064 4324
rect 2608 3836 2672 3840
rect 2608 3780 2612 3836
rect 2612 3780 2668 3836
rect 2668 3780 2672 3836
rect 2608 3776 2672 3780
rect 2688 3836 2752 3840
rect 2688 3780 2692 3836
rect 2692 3780 2748 3836
rect 2748 3780 2752 3836
rect 2688 3776 2752 3780
rect 2768 3836 2832 3840
rect 2768 3780 2772 3836
rect 2772 3780 2828 3836
rect 2828 3780 2832 3836
rect 2768 3776 2832 3780
rect 2848 3836 2912 3840
rect 2848 3780 2852 3836
rect 2852 3780 2908 3836
rect 2908 3780 2912 3836
rect 2848 3776 2912 3780
rect 4080 3836 4144 3840
rect 4080 3780 4084 3836
rect 4084 3780 4140 3836
rect 4140 3780 4144 3836
rect 4080 3776 4144 3780
rect 4160 3836 4224 3840
rect 4160 3780 4164 3836
rect 4164 3780 4220 3836
rect 4220 3780 4224 3836
rect 4160 3776 4224 3780
rect 4240 3836 4304 3840
rect 4240 3780 4244 3836
rect 4244 3780 4300 3836
rect 4300 3780 4304 3836
rect 4240 3776 4304 3780
rect 4320 3836 4384 3840
rect 4320 3780 4324 3836
rect 4324 3780 4380 3836
rect 4380 3780 4384 3836
rect 4320 3776 4384 3780
rect 5552 3836 5616 3840
rect 5552 3780 5556 3836
rect 5556 3780 5612 3836
rect 5612 3780 5616 3836
rect 5552 3776 5616 3780
rect 5632 3836 5696 3840
rect 5632 3780 5636 3836
rect 5636 3780 5692 3836
rect 5692 3780 5696 3836
rect 5632 3776 5696 3780
rect 5712 3836 5776 3840
rect 5712 3780 5716 3836
rect 5716 3780 5772 3836
rect 5772 3780 5776 3836
rect 5712 3776 5776 3780
rect 5792 3836 5856 3840
rect 5792 3780 5796 3836
rect 5796 3780 5852 3836
rect 5852 3780 5856 3836
rect 5792 3776 5856 3780
rect 7024 3836 7088 3840
rect 7024 3780 7028 3836
rect 7028 3780 7084 3836
rect 7084 3780 7088 3836
rect 7024 3776 7088 3780
rect 7104 3836 7168 3840
rect 7104 3780 7108 3836
rect 7108 3780 7164 3836
rect 7164 3780 7168 3836
rect 7104 3776 7168 3780
rect 7184 3836 7248 3840
rect 7184 3780 7188 3836
rect 7188 3780 7244 3836
rect 7244 3780 7248 3836
rect 7184 3776 7248 3780
rect 7264 3836 7328 3840
rect 7264 3780 7268 3836
rect 7268 3780 7324 3836
rect 7324 3780 7328 3836
rect 7264 3776 7328 3780
rect 3344 3292 3408 3296
rect 3344 3236 3348 3292
rect 3348 3236 3404 3292
rect 3404 3236 3408 3292
rect 3344 3232 3408 3236
rect 3424 3292 3488 3296
rect 3424 3236 3428 3292
rect 3428 3236 3484 3292
rect 3484 3236 3488 3292
rect 3424 3232 3488 3236
rect 3504 3292 3568 3296
rect 3504 3236 3508 3292
rect 3508 3236 3564 3292
rect 3564 3236 3568 3292
rect 3504 3232 3568 3236
rect 3584 3292 3648 3296
rect 3584 3236 3588 3292
rect 3588 3236 3644 3292
rect 3644 3236 3648 3292
rect 3584 3232 3648 3236
rect 4816 3292 4880 3296
rect 4816 3236 4820 3292
rect 4820 3236 4876 3292
rect 4876 3236 4880 3292
rect 4816 3232 4880 3236
rect 4896 3292 4960 3296
rect 4896 3236 4900 3292
rect 4900 3236 4956 3292
rect 4956 3236 4960 3292
rect 4896 3232 4960 3236
rect 4976 3292 5040 3296
rect 4976 3236 4980 3292
rect 4980 3236 5036 3292
rect 5036 3236 5040 3292
rect 4976 3232 5040 3236
rect 5056 3292 5120 3296
rect 5056 3236 5060 3292
rect 5060 3236 5116 3292
rect 5116 3236 5120 3292
rect 5056 3232 5120 3236
rect 6288 3292 6352 3296
rect 6288 3236 6292 3292
rect 6292 3236 6348 3292
rect 6348 3236 6352 3292
rect 6288 3232 6352 3236
rect 6368 3292 6432 3296
rect 6368 3236 6372 3292
rect 6372 3236 6428 3292
rect 6428 3236 6432 3292
rect 6368 3232 6432 3236
rect 6448 3292 6512 3296
rect 6448 3236 6452 3292
rect 6452 3236 6508 3292
rect 6508 3236 6512 3292
rect 6448 3232 6512 3236
rect 6528 3292 6592 3296
rect 6528 3236 6532 3292
rect 6532 3236 6588 3292
rect 6588 3236 6592 3292
rect 6528 3232 6592 3236
rect 7760 3292 7824 3296
rect 7760 3236 7764 3292
rect 7764 3236 7820 3292
rect 7820 3236 7824 3292
rect 7760 3232 7824 3236
rect 7840 3292 7904 3296
rect 7840 3236 7844 3292
rect 7844 3236 7900 3292
rect 7900 3236 7904 3292
rect 7840 3232 7904 3236
rect 7920 3292 7984 3296
rect 7920 3236 7924 3292
rect 7924 3236 7980 3292
rect 7980 3236 7984 3292
rect 7920 3232 7984 3236
rect 8000 3292 8064 3296
rect 8000 3236 8004 3292
rect 8004 3236 8060 3292
rect 8060 3236 8064 3292
rect 8000 3232 8064 3236
rect 2608 2748 2672 2752
rect 2608 2692 2612 2748
rect 2612 2692 2668 2748
rect 2668 2692 2672 2748
rect 2608 2688 2672 2692
rect 2688 2748 2752 2752
rect 2688 2692 2692 2748
rect 2692 2692 2748 2748
rect 2748 2692 2752 2748
rect 2688 2688 2752 2692
rect 2768 2748 2832 2752
rect 2768 2692 2772 2748
rect 2772 2692 2828 2748
rect 2828 2692 2832 2748
rect 2768 2688 2832 2692
rect 2848 2748 2912 2752
rect 2848 2692 2852 2748
rect 2852 2692 2908 2748
rect 2908 2692 2912 2748
rect 2848 2688 2912 2692
rect 4080 2748 4144 2752
rect 4080 2692 4084 2748
rect 4084 2692 4140 2748
rect 4140 2692 4144 2748
rect 4080 2688 4144 2692
rect 4160 2748 4224 2752
rect 4160 2692 4164 2748
rect 4164 2692 4220 2748
rect 4220 2692 4224 2748
rect 4160 2688 4224 2692
rect 4240 2748 4304 2752
rect 4240 2692 4244 2748
rect 4244 2692 4300 2748
rect 4300 2692 4304 2748
rect 4240 2688 4304 2692
rect 4320 2748 4384 2752
rect 4320 2692 4324 2748
rect 4324 2692 4380 2748
rect 4380 2692 4384 2748
rect 4320 2688 4384 2692
rect 5552 2748 5616 2752
rect 5552 2692 5556 2748
rect 5556 2692 5612 2748
rect 5612 2692 5616 2748
rect 5552 2688 5616 2692
rect 5632 2748 5696 2752
rect 5632 2692 5636 2748
rect 5636 2692 5692 2748
rect 5692 2692 5696 2748
rect 5632 2688 5696 2692
rect 5712 2748 5776 2752
rect 5712 2692 5716 2748
rect 5716 2692 5772 2748
rect 5772 2692 5776 2748
rect 5712 2688 5776 2692
rect 5792 2748 5856 2752
rect 5792 2692 5796 2748
rect 5796 2692 5852 2748
rect 5852 2692 5856 2748
rect 5792 2688 5856 2692
rect 7024 2748 7088 2752
rect 7024 2692 7028 2748
rect 7028 2692 7084 2748
rect 7084 2692 7088 2748
rect 7024 2688 7088 2692
rect 7104 2748 7168 2752
rect 7104 2692 7108 2748
rect 7108 2692 7164 2748
rect 7164 2692 7168 2748
rect 7104 2688 7168 2692
rect 7184 2748 7248 2752
rect 7184 2692 7188 2748
rect 7188 2692 7244 2748
rect 7244 2692 7248 2748
rect 7184 2688 7248 2692
rect 7264 2748 7328 2752
rect 7264 2692 7268 2748
rect 7268 2692 7324 2748
rect 7324 2692 7328 2748
rect 7264 2688 7328 2692
rect 3344 2204 3408 2208
rect 3344 2148 3348 2204
rect 3348 2148 3404 2204
rect 3404 2148 3408 2204
rect 3344 2144 3408 2148
rect 3424 2204 3488 2208
rect 3424 2148 3428 2204
rect 3428 2148 3484 2204
rect 3484 2148 3488 2204
rect 3424 2144 3488 2148
rect 3504 2204 3568 2208
rect 3504 2148 3508 2204
rect 3508 2148 3564 2204
rect 3564 2148 3568 2204
rect 3504 2144 3568 2148
rect 3584 2204 3648 2208
rect 3584 2148 3588 2204
rect 3588 2148 3644 2204
rect 3644 2148 3648 2204
rect 3584 2144 3648 2148
rect 4816 2204 4880 2208
rect 4816 2148 4820 2204
rect 4820 2148 4876 2204
rect 4876 2148 4880 2204
rect 4816 2144 4880 2148
rect 4896 2204 4960 2208
rect 4896 2148 4900 2204
rect 4900 2148 4956 2204
rect 4956 2148 4960 2204
rect 4896 2144 4960 2148
rect 4976 2204 5040 2208
rect 4976 2148 4980 2204
rect 4980 2148 5036 2204
rect 5036 2148 5040 2204
rect 4976 2144 5040 2148
rect 5056 2204 5120 2208
rect 5056 2148 5060 2204
rect 5060 2148 5116 2204
rect 5116 2148 5120 2204
rect 5056 2144 5120 2148
rect 6288 2204 6352 2208
rect 6288 2148 6292 2204
rect 6292 2148 6348 2204
rect 6348 2148 6352 2204
rect 6288 2144 6352 2148
rect 6368 2204 6432 2208
rect 6368 2148 6372 2204
rect 6372 2148 6428 2204
rect 6428 2148 6432 2204
rect 6368 2144 6432 2148
rect 6448 2204 6512 2208
rect 6448 2148 6452 2204
rect 6452 2148 6508 2204
rect 6508 2148 6512 2204
rect 6448 2144 6512 2148
rect 6528 2204 6592 2208
rect 6528 2148 6532 2204
rect 6532 2148 6588 2204
rect 6588 2148 6592 2204
rect 6528 2144 6592 2148
rect 7760 2204 7824 2208
rect 7760 2148 7764 2204
rect 7764 2148 7820 2204
rect 7820 2148 7824 2204
rect 7760 2144 7824 2148
rect 7840 2204 7904 2208
rect 7840 2148 7844 2204
rect 7844 2148 7900 2204
rect 7900 2148 7904 2204
rect 7840 2144 7904 2148
rect 7920 2204 7984 2208
rect 7920 2148 7924 2204
rect 7924 2148 7980 2204
rect 7980 2148 7984 2204
rect 7920 2144 7984 2148
rect 8000 2204 8064 2208
rect 8000 2148 8004 2204
rect 8004 2148 8060 2204
rect 8060 2148 8064 2204
rect 8000 2144 8064 2148
<< metal4 >>
rect 2600 7764 7336 8084
rect 2600 7104 2920 7764
rect 2600 7040 2608 7104
rect 2672 7040 2688 7104
rect 2752 7040 2768 7104
rect 2832 7040 2848 7104
rect 2912 7040 2920 7104
rect 2600 6016 2920 7040
rect 2600 5952 2608 6016
rect 2672 5952 2688 6016
rect 2752 5952 2768 6016
rect 2832 5952 2848 6016
rect 2912 5952 2920 6016
rect 2600 4928 2920 5952
rect 2600 4864 2608 4928
rect 2672 4864 2688 4928
rect 2752 4864 2768 4928
rect 2832 4864 2848 4928
rect 2912 4864 2920 4928
rect 2600 3840 2920 4864
rect 2600 3776 2608 3840
rect 2672 3776 2688 3840
rect 2752 3776 2768 3840
rect 2832 3776 2848 3840
rect 2912 3776 2920 3840
rect 2600 2752 2920 3776
rect 2600 2688 2608 2752
rect 2672 2688 2688 2752
rect 2752 2688 2768 2752
rect 2832 2688 2848 2752
rect 2912 2688 2920 2752
rect 2600 2128 2920 2688
rect 3336 7648 3656 7664
rect 3336 7584 3344 7648
rect 3408 7584 3424 7648
rect 3488 7584 3504 7648
rect 3568 7584 3584 7648
rect 3648 7584 3656 7648
rect 3336 6560 3656 7584
rect 3336 6496 3344 6560
rect 3408 6496 3424 6560
rect 3488 6496 3504 6560
rect 3568 6496 3584 6560
rect 3648 6496 3656 6560
rect 3336 5472 3656 6496
rect 3336 5408 3344 5472
rect 3408 5408 3424 5472
rect 3488 5408 3504 5472
rect 3568 5408 3584 5472
rect 3648 5408 3656 5472
rect 3336 4384 3656 5408
rect 3336 4320 3344 4384
rect 3408 4320 3424 4384
rect 3488 4320 3504 4384
rect 3568 4320 3584 4384
rect 3648 4320 3656 4384
rect 3336 3296 3656 4320
rect 3336 3232 3344 3296
rect 3408 3232 3424 3296
rect 3488 3232 3504 3296
rect 3568 3232 3584 3296
rect 3648 3232 3656 3296
rect 3336 2208 3656 3232
rect 3336 2144 3344 2208
rect 3408 2144 3424 2208
rect 3488 2144 3504 2208
rect 3568 2144 3584 2208
rect 3648 2144 3656 2208
rect 3336 1958 3656 2144
rect 4072 7104 4392 7764
rect 4072 7040 4080 7104
rect 4144 7040 4160 7104
rect 4224 7040 4240 7104
rect 4304 7040 4320 7104
rect 4384 7040 4392 7104
rect 4072 6016 4392 7040
rect 4072 5952 4080 6016
rect 4144 5952 4160 6016
rect 4224 5952 4240 6016
rect 4304 5952 4320 6016
rect 4384 5952 4392 6016
rect 4072 4928 4392 5952
rect 4072 4864 4080 4928
rect 4144 4864 4160 4928
rect 4224 4864 4240 4928
rect 4304 4864 4320 4928
rect 4384 4864 4392 4928
rect 4072 3840 4392 4864
rect 4072 3776 4080 3840
rect 4144 3776 4160 3840
rect 4224 3776 4240 3840
rect 4304 3776 4320 3840
rect 4384 3776 4392 3840
rect 4072 2752 4392 3776
rect 4072 2688 4080 2752
rect 4144 2688 4160 2752
rect 4224 2688 4240 2752
rect 4304 2688 4320 2752
rect 4384 2688 4392 2752
rect 4072 2128 4392 2688
rect 4808 7648 5128 7664
rect 4808 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5128 7648
rect 4808 6560 5128 7584
rect 4808 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5128 6560
rect 4808 5472 5128 6496
rect 4808 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5128 5472
rect 4808 4384 5128 5408
rect 4808 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5128 4384
rect 4808 3296 5128 4320
rect 4808 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5128 3296
rect 4808 2208 5128 3232
rect 4808 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5128 2208
rect 4808 1958 5128 2144
rect 5544 7104 5864 7764
rect 5544 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5864 7104
rect 5544 6016 5864 7040
rect 5544 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5864 6016
rect 5544 4928 5864 5952
rect 5544 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5864 4928
rect 5544 3840 5864 4864
rect 5544 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5864 3840
rect 5544 2752 5864 3776
rect 5544 2688 5552 2752
rect 5616 2688 5632 2752
rect 5696 2688 5712 2752
rect 5776 2688 5792 2752
rect 5856 2688 5864 2752
rect 5544 2128 5864 2688
rect 6280 7648 6600 7664
rect 6280 7584 6288 7648
rect 6352 7584 6368 7648
rect 6432 7584 6448 7648
rect 6512 7584 6528 7648
rect 6592 7584 6600 7648
rect 6280 6560 6600 7584
rect 6280 6496 6288 6560
rect 6352 6496 6368 6560
rect 6432 6496 6448 6560
rect 6512 6496 6528 6560
rect 6592 6496 6600 6560
rect 6280 5472 6600 6496
rect 6280 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6600 5472
rect 6280 4384 6600 5408
rect 6280 4320 6288 4384
rect 6352 4320 6368 4384
rect 6432 4320 6448 4384
rect 6512 4320 6528 4384
rect 6592 4320 6600 4384
rect 6280 3296 6600 4320
rect 6280 3232 6288 3296
rect 6352 3232 6368 3296
rect 6432 3232 6448 3296
rect 6512 3232 6528 3296
rect 6592 3232 6600 3296
rect 6280 2208 6600 3232
rect 6280 2144 6288 2208
rect 6352 2144 6368 2208
rect 6432 2144 6448 2208
rect 6512 2144 6528 2208
rect 6592 2144 6600 2208
rect 6280 1958 6600 2144
rect 7016 7104 7336 7764
rect 7016 7040 7024 7104
rect 7088 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7336 7104
rect 7016 6016 7336 7040
rect 7016 5952 7024 6016
rect 7088 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7336 6016
rect 7016 4928 7336 5952
rect 7016 4864 7024 4928
rect 7088 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7336 4928
rect 7016 3840 7336 4864
rect 7016 3776 7024 3840
rect 7088 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7336 3840
rect 7016 2752 7336 3776
rect 7016 2688 7024 2752
rect 7088 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7336 2752
rect 7016 2128 7336 2688
rect 7752 7648 8072 7664
rect 7752 7584 7760 7648
rect 7824 7584 7840 7648
rect 7904 7584 7920 7648
rect 7984 7584 8000 7648
rect 8064 7584 8072 7648
rect 7752 6560 8072 7584
rect 7752 6496 7760 6560
rect 7824 6496 7840 6560
rect 7904 6496 7920 6560
rect 7984 6496 8000 6560
rect 8064 6496 8072 6560
rect 7752 5472 8072 6496
rect 7752 5408 7760 5472
rect 7824 5408 7840 5472
rect 7904 5408 7920 5472
rect 7984 5408 8000 5472
rect 8064 5408 8072 5472
rect 7752 4384 8072 5408
rect 7752 4320 7760 4384
rect 7824 4320 7840 4384
rect 7904 4320 7920 4384
rect 7984 4320 8000 4384
rect 8064 4320 8072 4384
rect 7752 3296 8072 4320
rect 7752 3232 7760 3296
rect 7824 3232 7840 3296
rect 7904 3232 7920 3296
rect 7984 3232 8000 3296
rect 8064 3232 8072 3296
rect 7752 2208 8072 3232
rect 7752 2144 7760 2208
rect 7824 2144 7840 2208
rect 7904 2144 7920 2208
rect 7984 2144 8000 2208
rect 8064 2144 8072 2208
rect 7752 1958 8072 2144
rect 3336 1638 8072 1958
use sky130_fd_sc_hd__clkbuf_2  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _12_
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _13_
timestamp 1704896540
transform 1 0 4140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2760 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _16_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1704896540
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _20_
timestamp 1704896540
transform 1 0 2576 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _21_
timestamp 1704896540
transform 1 0 3404 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1704896540
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2852 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1704896540
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _26_
timestamp 1704896540
transform 1 0 2576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _27_
timestamp 1704896540
transform 1 0 4140 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1704896540
transform -1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _29_
timestamp 1704896540
transform -1 0 4324 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1704896540
transform -1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _31_
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _32_
timestamp 1704896540
transform -1 0 3680 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1704896540
transform 1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _34_
timestamp 1704896540
transform 1 0 5244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1704896540
transform 1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48
timestamp 1704896540
transform 1 0 6440 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7268 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_13
timestamp 1704896540
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_25
timestamp 1704896540
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_37
timestamp 1704896540
transform 1 0 5428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1704896540
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_22
timestamp 1704896540
transform 1 0 4048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1704896540
transform 1 0 6900 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_3
timestamp 1704896540
transform 1 0 2300 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_19
timestamp 1704896540
transform 1 0 3772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_25
timestamp 1704896540
transform 1 0 4324 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_30
timestamp 1704896540
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_42
timestamp 1704896540
transform 1 0 5888 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1704896540
transform 1 0 6992 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1704896540
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1704896540
transform 1 0 2852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1704896540
transform 1 0 3956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1704896540
transform 1 0 6900 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 1704896540
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_20
timestamp 1704896540
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_32
timestamp 1704896540
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_44
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1704896540
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_9
timestamp 1704896540
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1704896540
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_35
timestamp 1704896540
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_47
timestamp 1704896540
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_59
timestamp 1704896540
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_22
timestamp 1704896540
transform 1 0 4048 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_30
timestamp 1704896540
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_34
timestamp 1704896540
transform 1 0 5152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_47
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1704896540
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1704896540
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_34
timestamp 1704896540
transform 1 0 5152 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_42
timestamp 1704896540
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_54
timestamp 1704896540
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1704896540
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_35
timestamp 1704896540
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1704896540
transform 1 0 7268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1704896540
transform -1 0 4324 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1704896540
transform -1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1704896540
transform -1 0 5244 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1704896540
transform 1 0 5520 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1704896540
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1704896540
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1704896540
transform 1 0 6072 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1704896540
transform 1 0 2852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1704896540
transform -1 0 2852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1704896540
transform -1 0 2852 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1704896540
transform -1 0 2852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1704896540
transform -1 0 2852 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1704896540
transform -1 0 3956 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1704896540
transform -1 0 2852 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1704896540
transform -1 0 2852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 1704896540
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 1704896540
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 1704896540
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 1704896540
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 1704896540
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 1704896540
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 1704896540
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 1704896540
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 1704896540
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 1704896540
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 1704896540
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 1704896540
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 1704896540
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 1704896540
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 1704896540
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 1704896540
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 1704896540
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 1704896540
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 1704896540
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 1704896540
transform 1 0 4600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 1704896540
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string GDS_END 213802
string GDS_FILE ../gds/decoder_p.gds
string GDS_START 81952
<< end >>
