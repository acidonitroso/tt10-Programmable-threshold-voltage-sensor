VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decoder_p
  CLASS BLOCK ;
  FOREIGN decoder_p ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 50.000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 38.760 10.640 40.360 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.400 10.640 33.000 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.040 10.640 25.640 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.680 10.640 18.280 38.320 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 35.080 10.640 36.680 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.720 10.640 29.320 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.360 10.640 21.960 38.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.000 10.640 14.600 38.320 ;
    END
  END VPWR
  PIN in[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 2.000 ;
    END
  END in[0]
  PIN in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.000 ;
    END
  END in[1]
  PIN in[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.000 ;
    END
  END in[2]
  PIN n_d[0]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.770 48.000 4.050 50.000 ;
    END
  END n_d[0]
  PIN n_d[1]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 48.000 10.030 50.000 ;
    END
  END n_d[1]
  PIN n_d[2]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 15.730 48.000 16.010 50.000 ;
    END
  END n_d[2]
  PIN n_d[3]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 21.710 48.000 21.990 50.000 ;
    END
  END n_d[3]
  PIN n_d[4]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 27.690 48.000 27.970 50.000 ;
    END
  END n_d[4]
  PIN n_d[5]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 33.670 48.000 33.950 50.000 ;
    END
  END n_d[5]
  PIN n_d[6]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 39.650 48.000 39.930 50.000 ;
    END
  END n_d[6]
  PIN n_d[7]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.630 48.000 45.910 50.000 ;
    END
  END n_d[7]
  PIN y_d[0]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 2.000 6.080 ;
    END
  END y_d[0]
  PIN y_d[1]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END y_d[1]
  PIN y_d[2]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.000 16.960 ;
    END
  END y_d[2]
  PIN y_d[3]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.000 22.400 ;
    END
  END y_d[3]
  PIN y_d[4]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 2.000 27.840 ;
    END
  END y_d[4]
  PIN y_d[5]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.000 33.280 ;
    END
  END y_d[5]
  PIN y_d[6]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.000 38.720 ;
    END
  END y_d[6]
  PIN y_d[7]
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.000 44.160 ;
    END
  END y_d[7]
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 39.560 38.165 ;
      LAYER met1 ;
        RECT 3.750 10.640 45.930 38.320 ;
      LAYER met2 ;
        RECT 4.330 47.720 9.470 48.690 ;
        RECT 10.310 47.720 15.450 48.690 ;
        RECT 16.290 47.720 21.430 48.690 ;
        RECT 22.270 47.720 27.410 48.690 ;
        RECT 28.250 47.720 33.390 48.690 ;
        RECT 34.230 47.720 39.370 48.690 ;
        RECT 40.210 47.720 45.350 48.690 ;
        RECT 3.780 2.280 45.900 47.720 ;
        RECT 3.780 2.000 8.090 2.280 ;
        RECT 8.930 2.000 24.650 2.280 ;
        RECT 25.490 2.000 41.210 2.280 ;
        RECT 42.050 2.000 45.900 2.280 ;
      LAYER met3 ;
        RECT 2.400 43.160 40.350 44.025 ;
        RECT 2.000 39.120 40.350 43.160 ;
        RECT 2.400 37.720 40.350 39.120 ;
        RECT 2.000 33.680 40.350 37.720 ;
        RECT 2.400 32.280 40.350 33.680 ;
        RECT 2.000 28.240 40.350 32.280 ;
        RECT 2.400 26.840 40.350 28.240 ;
        RECT 2.000 22.800 40.350 26.840 ;
        RECT 2.400 21.400 40.350 22.800 ;
        RECT 2.000 17.360 40.350 21.400 ;
        RECT 2.400 15.960 40.350 17.360 ;
        RECT 2.000 11.920 40.350 15.960 ;
        RECT 2.400 10.520 40.350 11.920 ;
        RECT 2.000 6.480 40.350 10.520 ;
        RECT 2.400 5.615 40.350 6.480 ;
      LAYER met4 ;
        RECT 13.000 38.720 40.360 40.420 ;
        RECT 15.000 10.240 16.280 38.720 ;
        RECT 18.680 10.240 19.960 38.720 ;
        RECT 22.360 10.240 23.640 38.720 ;
        RECT 26.040 10.240 27.320 38.720 ;
        RECT 29.720 10.240 31.000 38.720 ;
        RECT 33.400 10.240 34.680 38.720 ;
        RECT 37.080 10.240 38.360 38.720 ;
        RECT 13.000 8.190 40.360 10.240 ;
  END
END decoder_p
END LIBRARY

