magic
tech sky130A
magscale 1 2
timestamp 1750694016
<< viali >>
rect 252 4498 340 4692
rect 764 4502 852 4696
<< metal1 >>
rect 62 7112 1034 7574
rect 226 4696 870 4704
rect 226 4692 764 4696
rect 226 4498 252 4692
rect 340 4502 764 4692
rect 852 4502 870 4696
rect 340 4498 870 4502
rect 226 4488 870 4498
rect 498 4006 702 4488
rect 786 4006 1090 4220
rect 498 3802 1090 4006
rect 786 3616 1090 3802
rect 786 3306 1090 3312
rect -447 1721 -225 1727
rect -447 1160 -225 1499
rect -458 530 308 1160
<< via1 >>
rect 786 3312 1090 3616
rect -447 1499 -225 1721
<< metal2 >>
rect 780 3312 786 3616
rect 1090 3312 1096 3616
rect 786 3091 1090 3100
rect -447 2065 -225 2074
rect -447 1721 -225 1843
rect -453 1499 -447 1721
rect -225 1499 -219 1721
<< via2 >>
rect 786 3312 1090 3404
rect 786 3100 1090 3312
rect -447 1843 -225 2065
<< metal3 >>
rect 781 3404 1095 3409
rect 781 3095 786 3404
rect 1090 3095 1095 3404
rect 786 2882 1090 2888
rect -447 2385 -225 2391
rect -447 2070 -225 2163
rect -452 2065 -220 2070
rect -452 1843 -447 2065
rect -225 1843 -220 2065
rect -452 1838 -220 1843
<< via3 >>
rect 786 3100 1090 3192
rect 786 2888 1090 3100
rect -447 2163 -225 2385
<< metal4 >>
rect -447 2386 -225 7711
rect 785 3192 1091 3193
rect 785 2888 786 3192
rect 1090 2888 1091 3192
rect 785 2887 1091 2888
rect 786 2720 1090 2887
rect -448 2385 -224 2386
rect -448 2163 -447 2385
rect -225 2163 -224 2385
rect -448 2162 -224 2163
use sky130_fd_pr__res_high_po_0p35_M898NC  XR9
timestamp 1749663830
transform 1 0 148 0 1 4139
box -201 -3592 201 3592
use sky130_fd_pr__res_high_po_0p35_J32JWA  XR10
timestamp 1749663830
transform 1 0 953 0 1 5678
box -201 -2052 201 2052
<< end >>
