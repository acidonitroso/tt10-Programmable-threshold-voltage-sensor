magic
tech sky130A
magscale 1 2
timestamp 1750694058
<< viali >>
rect -454 4798 -406 5002
rect 128 4800 180 5000
<< metal1 >>
rect -638 7078 388 7520
rect -474 5002 206 5014
rect -474 4798 -454 5002
rect -406 5000 206 5002
rect -406 4800 128 5000
rect 180 4800 206 5000
rect -406 4798 206 4800
rect -474 4774 206 4798
rect -1098 3054 -878 3060
rect -1098 2488 -878 2834
rect -1098 2478 -486 2488
rect -1098 2072 -474 2478
rect -1098 2068 -878 2072
rect -694 2068 -474 2072
rect -204 1004 -4 4774
rect 138 1004 474 1090
rect -204 804 474 1004
rect 138 632 474 804
rect 138 290 474 296
<< via1 >>
rect -1098 2834 -878 3054
rect 138 296 474 632
<< metal2 >>
rect -1098 3334 -878 3343
rect -1098 3054 -878 3114
rect -1104 2834 -1098 3054
rect -878 2834 -872 3054
rect 132 296 138 632
rect 474 296 480 632
rect 138 284 474 296
rect 138 -61 474 -52
<< via2 >>
rect -1098 3114 -878 3334
rect 138 -52 474 284
<< metal3 >>
rect -1098 3700 -878 3706
rect -1098 3339 -878 3480
rect -1103 3334 -873 3339
rect -1103 3114 -1098 3334
rect -878 3114 -873 3334
rect -1103 3109 -873 3114
rect 133 284 479 289
rect 133 -52 138 284
rect 474 -52 479 284
rect 133 -57 479 -52
rect 138 -60 474 -57
rect 138 -402 474 -396
<< via3 >>
rect -1098 3480 -878 3700
rect 138 -396 474 -60
<< metal4 >>
rect -1098 3701 -878 7902
rect -1099 3700 -877 3701
rect -1099 3480 -1098 3700
rect -878 3480 -877 3700
rect -1099 3479 -877 3480
rect 137 -60 475 -59
rect 137 -396 138 -60
rect 474 -396 475 -60
rect 137 -397 475 -396
rect 138 -600 474 -397
use sky130_fd_pr__res_high_po_0p35_A5V4E5  XR1
timestamp 1749662202
transform 1 0 -581 0 1 4792
box -201 -2892 201 2892
use sky130_fd_pr__res_high_po_0p35_M898NC  XR4
timestamp 1749663830
transform 1 0 301 0 1 4098
box -201 -3592 201 3592
<< end >>
