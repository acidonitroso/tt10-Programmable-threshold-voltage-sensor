* NGSPICE file created from decoder_p_parax.ext - technology: sky130A

.subckt decoder_p n_d[1] n_d[3] n_d[4] n_d[6] y_d[0] y_d[1] y_d[2] y_d[3] y_d[4] y_d[5] y_d[6] y_d[7] in[0] in[2] n_d[5] n_d[0] in[1] n_d[2] n_d[7] VGND VPWR
X0 VPWR.t256 VGND.t504 VPWR.t255 VPWR.t254 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 _01_.t1 a_3707_3311# VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X2 VGND.t66 a_3571_4074# net15 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3 a_3307_7379# net6 VGND.t356 VGND.t355 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4 n_d[0].t7 a_2939_6549# VGND.t236 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND.t360 a_3019_7338# net18 VGND.t359 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X6 VGND.t208 a_3755_5639# _08_ VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR.t276 a_2879_2223# y_d[0].t3 VPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X8 VPWR.t61 a_5137_2388# net2 VPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X9 _10_ a_3155_5056# VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X10 a_4031_6740# _05_ VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X11 VGND.t302 a_2387_7379# y_d[6].t7 VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 n_d[1].t7 a_3859_7379# VGND.t354 VGND.t353 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X13 a_3373_3561# _02_ a_3289_3561# VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR.t321 a_6099_7119# n_d[7].t3 VPWR.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X15 a_4509_6147# net2 a_4437_6147# VPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 VPWR.t253 VGND.t505 VPWR.t252 VPWR.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X17 a_4399_7338# _04_ VPWR.t379 VPWR.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X18 VGND.t346 VPWR.t491 VGND.t345 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X19 VPWR.t397 _02_ a_3155_5056# VPWR.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X20 VGND.t404 _02_ a_5849_6147# VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X21 VGND.t286 a_4443_3855# _00_ VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_3148_4215# a_2961_3855# a_3061_3971# VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X23 VGND.t227 a_2879_2223# y_d[0].t7 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 _05_ a_3619_6147# VGND.t461 VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X25 VGND.t435 a_2869_6147# a_2975_6147# VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 n_d[7].t2 a_6099_7119# VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X27 VGND.t469 a_2387_6549# y_d[7].t7 VGND.t468 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VPWR.t329 a_2387_7379# y_d[6].t3 VPWR.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR.t360 net9 a_6651_7119# VPWR.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X30 VPWR.t250 VGND.t506 VPWR.t249 VPWR.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X31 y_d[4].t3 a_2387_5461# VPWR.t420 VPWR.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 a_2939_6549# net4 VPWR.t434 VPWR.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X33 VPWR.t248 VGND.t507 VPWR.t247 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X34 VPWR.t373 net1 a_4509_6147# VPWR.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X35 VPWR.t438 a_2387_3027# y_d[2].t3 VPWR.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X36 VPWR.t246 VGND.t508 VPWR.t245 VPWR.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X37 VGND.t235 a_2939_6549# n_d[0].t6 VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 VPWR.t266 a_3491_6549# y_d[5].t3 VPWR.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X39 a_3309_5309# _01_.t4 a_3237_5309# VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X40 net1 a_3431_2223# VPWR.t258 VPWR.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X41 VGND.t94 VPWR.t492 VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X42 VPWR.t55 _01_.t5 a_5297_6147# VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X43 VGND.t97 VPWR.t493 VGND.t96 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X44 VGND.t191 VPWR.t494 VGND.t190 VGND.t189 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X45 n_d[4].t3 a_5547_7119# VPWR.t469 VPWR.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X46 VPWR.t243 VGND.t509 VPWR.t242 VPWR.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X47 y_d[2].t2 a_2387_3027# VPWR.t437 VPWR.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X48 y_d[5].t2 a_3491_6549# VPWR.t264 VPWR.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X49 VPWR.t240 VGND.t510 VPWR.t239 VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X50 VGND.t133 a_5137_2388# net2 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X51 a_5008_5487# _01_.t6 a_4924_5487# VGND.t249 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 a_3061_3971# net1 VPWR.t371 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X53 a_4031_6740# _05_ VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X54 VGND.t352 a_3859_7379# n_d[1].t6 VGND.t351 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X55 VPWR.t238 VGND.t511 VPWR.t237 VPWR.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X56 a_3057_6147# a_2869_6147# a_2975_6147# VPWR.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X57 net11 _00_ VPWR.t489 VPWR.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X58 VPWR.t412 a_7437_2388# net3 VPWR.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X59 VGND.t501 _00_ a_4745_5533# VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X60 a_2667_3463# _02_ VGND.t402 VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X61 a_2387_2197# net13 VPWR.t457 VPWR.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X62 a_2667_3463# _02_ VPWR.t395 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X63 a_3755_5639# a_4028_5467# a_3986_5493# VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X64 VPWR.t235 VGND.t512 VPWR.t234 VPWR.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X65 a_3491_6549# net17 VGND.t455 VGND.t454 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X66 VGND.t194 VPWR.t495 VGND.t193 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X67 VGND.t178 net8 a_5547_7119# VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X68 VGND.t128 VPWR.t496 VGND.t127 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X69 net7 a_4745_5533# VPWR.t53 VPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X70 VPWR.t428 a_5687_6740# net19 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X71 VPWR.t317 a_6099_7119# n_d[7].t1 VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X72 VGND.t131 VPWR.t497 VGND.t130 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X73 VPWR.t286 a_2939_6549# n_d[0].t3 VPWR.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X74 VPWR.t232 VGND.t513 VPWR.t231 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X75 y_d[6].t2 a_2387_7379# VPWR.t327 VPWR.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X76 VGND.t264 VPWR.t498 VGND.t263 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X77 VPWR.t350 a_3859_7379# n_d[1].t3 VPWR.t349 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X78 VPWR.t302 _01_.t7 a_3384_5467# VPWR.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X79 VGND.t267 VPWR.t499 VGND.t266 VGND.t265 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X80 VPWR.t93 a_6651_7119# n_d[5].t3 VPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X81 VPWR.t229 VGND.t514 VPWR.t228 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X82 VPWR.t227 VGND.t515 VPWR.t226 VPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X83 VGND.t341 VPWR.t500 VGND.t340 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X84 a_3859_7379# net5 VPWR.t402 VPWR.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X85 net1 a_3431_2223# VGND.t210 VGND.t209 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X86 a_2821_3561# _01_.t8 a_2737_3561# VPWR.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X87 VGND.t314 _01_.t9 net16 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X88 VPWR.t37 net3 a_4443_3855# VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X89 VPWR.t422 a_3111_5639# _09_ VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X90 VPWR.t467 a_5547_7119# n_d[4].t2 VPWR.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X91 VPWR.t456 a_2387_6549# y_d[7].t3 VPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X92 VPWR.t436 a_2387_3027# y_d[2].t1 VPWR.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X93 VPWR.t224 VGND.t516 VPWR.t223 VPWR.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X94 VPWR.t487 _00_ a_3045_2767# VPWR.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X95 a_2821_4943# _02_ a_2737_4943# VPWR.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X96 VGND.t418 a_7437_2388# net3 VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X97 net10 _00_ VPWR.t485 VPWR.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X98 n_d[4].t1 a_5547_7119# VPWR.t465 VPWR.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X99 y_d[7].t2 a_2387_6549# VPWR.t455 VPWR.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X100 VGND.t70 a_4167_3311# _02_ VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 _06_ a_3061_3971# VGND.t475 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X102 a_2387_5461# net16 VGND.t358 VGND.t357 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X103 _00_ a_4443_3855# VPWR.t313 VPWR.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X104 a_3111_5639# net3 VPWR.t35 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X105 a_2961_3855# _00_ VPWR.t483 VPWR.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X106 a_3261_5493# net3 VGND.t46 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X107 VGND.t433 a_5687_6740# net19 VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X108 VPWR.t221 VGND.t517 VPWR.t220 VPWR.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X109 n_d[7].t0 a_6099_7119# VPWR.t315 VPWR.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X110 n_d[0].t2 a_2939_6549# VPWR.t284 VPWR.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X111 VGND.t147 net12 a_2879_2223# VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X112 VPWR.t369 net1 a_3707_3311# VPWR.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X113 VPWR.t219 VGND.t518 VPWR.t218 VPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X114 VGND.t344 VPWR.t501 VGND.t343 VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X115 VPWR.t358 a_4399_7338# net5 VPWR.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X116 VGND.t400 _02_ a_4028_5467# VGND.t399 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X117 VGND.t44 net3 a_2975_6147# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X118 net7 _02_ VPWR.t392 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X119 VGND.t259 VPWR.t502 VGND.t258 VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X120 VGND.t108 net11 a_6099_7119# VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X121 net12 _01_.t10 VGND.t272 VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X122 n_d[2].t7 a_3307_7379# VGND.t143 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X123 VGND.t378 net1 a_2376_6263# VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X124 VPWR.t217 VGND.t519 VPWR.t216 VPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X125 y_d[2].t0 a_2387_3027# VPWR.t435 VPWR.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X126 a_3019_7338# _09_ VPWR.t85 VPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X127 VGND.t274 _01_.t11 a_5297_6147# VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X128 net17 a_3615_4943# VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X129 VPWR.t463 a_5547_7119# n_d[4].t0 VPWR.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X130 VPWR.t454 a_2387_6549# y_d[7].t1 VPWR.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X131 VPWR.t444 a_2376_6263# _03_ VPWR.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X132 VPWR.t215 VGND.t520 VPWR.t214 VPWR.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X133 n_d[2].t3 a_3307_7379# VPWR.t71 VPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X134 VPWR.t212 VGND.t521 VPWR.t211 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X135 _01_.t3 a_3707_3311# VGND.t64 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X136 VPWR.t282 a_2939_6549# n_d[0].t1 VPWR.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X137 n_d[5].t7 a_6651_7119# VGND.t204 VGND.t203 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X138 a_3307_7379# net6 VPWR.t352 VPWR.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X139 VGND.t42 net3 a_3619_6147# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 y_d[3].t7 a_2387_4373# VGND.t416 VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X141 a_3342_5493# net2 a_3261_5493# VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X142 net13 _02_ VGND.t398 VGND.t397 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X143 VGND.t261 VPWR.t503 VGND.t260 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X144 a_2737_3561# a_2667_3463# net14 VPWR.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X145 a_4249_6147# net3 VPWR.t33 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X146 _02_ a_4167_3311# VPWR.t51 VPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X147 n_d[1].t2 a_3859_7379# VPWR.t348 VPWR.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X148 VGND.t50 VPWR.t504 VGND.t49 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X149 VPWR.t333 _01_.t12 net11 VPWR.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X150 VPWR.t22 net2 a_3111_5639# VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X151 VPWR.t43 a_3707_3311# _01_.t0 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X152 VPWR.t298 a_2387_2197# y_d[1].t3 VPWR.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X153 net17 a_3615_4943# VGND.t100 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X154 a_2737_4943# a_2667_5175# net16 VPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X155 VGND.t350 a_3859_7379# n_d[1].t5 VGND.t349 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X156 VPWR.t209 VGND.t522 VPWR.t208 VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X157 net10 a_5297_6147# a_5560_6351# VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X158 VPWR.t342 a_7111_6575# n_d[6].t3 VPWR.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X159 VPWR.t432 a_4307_6740# net4 VPWR.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X160 VPWR.t207 VGND.t523 VPWR.t206 VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X161 y_d[7].t0 a_2387_6549# VPWR.t453 VPWR.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X162 y_d[1].t2 a_2387_2197# VPWR.t296 VPWR.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X163 VPWR.t481 _00_ a_3373_3561# VPWR.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X164 VPWR.t205 VGND.t524 VPWR.t204 VPWR.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X165 a_3513_6147# net2 VPWR.t20 VPWR.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X166 VGND.t202 a_6651_7119# n_d[5].t6 VGND.t201 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X167 VGND.t52 VPWR.t505 VGND.t51 VGND.t48 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X168 a_4399_7338# _04_ VGND.t384 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X169 a_2387_3027# net14 VGND.t382 VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X170 _10_ a_3155_5056# VPWR.t12 VPWR.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X171 VGND.t380 net10 a_7111_6575# VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X172 VPWR.t202 VGND.t525 VPWR.t201 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X173 VGND.t57 VPWR.t506 VGND.t56 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X174 a_5560_6351# _02_ a_5476_6351# VGND.t396 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 VPWR.t346 a_3859_7379# n_d[1].t1 VPWR.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X176 a_2387_4373# net15 VPWR.t83 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X177 _04_ a_2975_6147# VPWR.t426 VPWR.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X178 VGND.t414 a_2387_4373# y_d[3].t6 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X179 n_d[2].t6 a_3307_7379# VGND.t141 VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X180 VGND.t60 VPWR.t507 VGND.t59 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X181 a_2387_2197# net13 VGND.t471 VGND.t470 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X182 VGND.t14 VPWR.t508 VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X183 y_d[3].t5 a_2387_4373# VGND.t412 VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X184 a_2667_5175# _00_ VPWR.t479 VPWR.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X185 VPWR.t199 VGND.t526 VPWR.t198 VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X186 VGND.t17 VPWR.t509 VGND.t16 VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X187 VPWR.t79 net8 a_5547_7119# VPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X188 a_4779_7379# net7 VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X189 VPWR.t196 VGND.t527 VPWR.t195 VPWR.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X190 VGND.t122 VPWR.t510 VGND.t121 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X191 VGND.t439 a_4307_6740# net4 VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X192 VPWR.t193 VGND.t528 VPWR.t192 VPWR.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X193 VPWR.t190 VGND.t529 VPWR.t189 VPWR.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X194 a_3289_3561# a_3219_3463# net13 VPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X195 VPWR.t294 a_2387_2197# y_d[1].t1 VPWR.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X196 a_4355_6147# net2 VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X197 a_3571_4074# _06_ VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X198 VPWR.t187 VGND.t530 VPWR.t186 VPWR.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X199 a_2869_6147# net1 VPWR.t367 VPWR.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X200 a_5687_6740# _10_ VPWR.t278 VPWR.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X201 n_d[5].t5 a_6651_7119# VGND.t200 VGND.t199 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X202 VPWR.t340 a_7111_6575# n_d[6].t2 VPWR.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X203 a_2387_7379# net18 VGND.t238 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X204 net14 _01_.t13 VGND.t312 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X205 _05_ a_3619_6147# VPWR.t452 VPWR.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X206 VPWR.t400 a_4031_6740# net6 VPWR.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X207 VGND.t125 VPWR.t511 VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X208 net9 a_5849_6147# a_6112_6351# VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X209 VGND.t305 VPWR.t512 VGND.t304 VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X210 VPWR.t184 VGND.t531 VPWR.t183 VPWR.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X211 VPWR.t181 VGND.t532 VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X212 VGND.t139 a_3307_7379# n_d[2].t5 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X213 VGND.t395 _02_ a_3309_5309# VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X214 a_2387_6549# net19 VGND.t366 VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X215 VPWR.t18 net2 a_3061_3971# VPWR.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X216 a_2607_6147# net1 a_2511_6147# VPWR.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X217 VGND.t294 a_6099_7119# n_d[7].t7 VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X218 VGND.t308 VPWR.t513 VGND.t307 VGND.t306 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X219 VPWR.t97 a_3755_5639# _08_ VPWR.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X220 VPWR.t477 _00_ a_2821_3561# VPWR.t476 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X221 VGND.t410 a_2387_4373# y_d[3].t4 VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X222 a_6112_6351# _01_.t14 a_6028_6351# VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 a_4249_6147# net3 VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X224 VPWR.t178 VGND.t533 VPWR.t177 VPWR.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X225 VPWR.t176 VGND.t534 VPWR.t175 VPWR.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X226 a_3129_6147# net2 a_3057_6147# VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X227 VPWR.t173 VGND.t535 VPWR.t172 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X228 n_d[0].t5 a_2939_6549# VGND.t233 VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X229 VGND.t88 VPWR.t514 VGND.t87 VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X230 n_d[7].t6 a_6099_7119# VGND.t292 VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X231 VGND.t91 VPWR.t515 VGND.t90 VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X232 VGND.t376 net1 a_3707_3311# VGND.t375 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X233 VPWR.t75 in[0].t0 a_3431_2223# VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X234 VPWR.t308 _01_.t15 a_2821_4943# VPWR.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X235 VPWR.t69 a_3307_7379# n_d[2].t2 VPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X236 y_d[1].t0 a_2387_2197# VPWR.t292 VPWR.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X237 VPWR.t424 a_2961_3855# a_3061_3971# VPWR.t423 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X238 _07_ a_4355_6147# VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X239 a_5687_6740# _10_ VGND.t229 VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X240 n_d[1].t4 a_3859_7379# VGND.t348 VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X241 a_3755_5639# net3 VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X242 a_5353_6575# _02_ VGND.t393 VGND.t392 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X243 n_d[6].t1 a_7111_6575# VPWR.t338 VPWR.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X244 VPWR.t171 VGND.t536 VPWR.t170 VPWR.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X245 VGND.t406 a_4031_6740# net6 VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X246 VPWR.t311 a_4443_3855# _00_ VPWR.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X247 a_3905_5493# net3 VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X248 VPWR.t59 net11 a_6099_7119# VPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X249 VPWR.t168 VGND.t537 VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X250 VPWR.t29 net3 a_3129_6147# VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X251 VGND.t167 VPWR.t516 VGND.t166 VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X252 a_3513_6147# net2 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X253 n_d[4].t7 a_5547_7119# VGND.t483 VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X254 VPWR.t15 net2 a_4167_3311# VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X255 _06_ a_3061_3971# VPWR.t461 VPWR.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X256 VGND.t362 a_4399_7338# net5 VGND.t361 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X257 VPWR.t390 _02_ a_4028_5467# VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X258 n_d[1].t0 a_3859_7379# VPWR.t344 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X259 a_3571_4074# _06_ VGND.t459 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X260 a_6028_6351# _00_ VGND.t499 VGND.t498 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X261 VPWR.t165 VGND.t538 VPWR.t164 VPWR.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X262 VPWR.t441 _01_.t16 net7 VPWR.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X263 VPWR.t162 VGND.t539 VPWR.t161 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X264 VGND.t391 _02_ net12 VGND.t390 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X265 VGND.t170 VPWR.t517 VGND.t169 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X266 net8 a_4903_6575# VPWR.t459 VPWR.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X267 VGND.t137 a_3307_7379# n_d[2].t4 VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X268 n_d[3].t7 a_4779_7379# VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X269 a_3755_5639# a_4028_5467# VPWR.t290 VPWR.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X270 a_2376_6263# net2 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X271 VGND.t82 VPWR.t518 VGND.t81 VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X272 a_3019_7338# _09_ VGND.t196 VGND.t195 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X273 VGND.t290 a_6099_7119# n_d[7].t5 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X274 a_5137_2388# in[1].t0 VPWR.t304 VPWR.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X275 VPWR.t159 VGND.t540 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X276 VGND.t72 in[0].t1 a_3431_2223# VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X277 VGND.t85 VPWR.t519 VGND.t84 VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X278 VGND.t503 a_4249_6147# a_4355_6147# VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X279 a_3045_2767# _01_.t17 a_2961_2767# VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 y_d[4].t7 a_2387_5461# VGND.t426 VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X281 a_3491_6549# net17 VPWR.t446 VPWR.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X282 VGND.t149 VPWR.t520 VGND.t148 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X283 a_2939_6549# net4 VGND.t441 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X284 VGND.t218 a_3491_6549# y_d[5].t7 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X285 VGND.t198 a_6651_7119# n_d[5].t4 VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X286 VPWR.t410 a_2387_4373# y_d[3].t3 VPWR.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X287 VGND.t437 a_2667_3463# net14 VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X288 VGND.t152 VPWR.t521 VGND.t151 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X289 VPWR.t27 net3 a_3773_6147# VPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X290 _02_ a_4167_3311# VGND.t68 VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X291 VPWR.t67 a_3307_7379# n_d[2].t1 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X292 VGND.t62 a_3707_3311# _01_.t2 VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X293 a_2869_6147# net1 VGND.t374 VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X294 VGND.t339 a_7111_6575# n_d[6].t7 VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X295 VGND.t481 a_5547_7119# n_d[4].t6 VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X296 y_d[3].t2 a_2387_4373# VPWR.t408 VPWR.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X297 VGND.t161 VPWR.t522 VGND.t160 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X298 n_d[6].t0 a_7111_6575# VPWR.t336 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X299 a_2376_6263# net2 a_2607_6147# VPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X300 VGND.t164 VPWR.t523 VGND.t163 VGND.t162 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X301 a_3986_5493# net1 a_3905_5493# VGND.t372 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X302 net11 _00_ a_5437_6575# VGND.t497 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X303 VGND.t451 a_3513_6147# a_3619_6147# VGND.t450 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X304 VPWR.t156 VGND.t541 VPWR.t155 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X305 a_4437_6147# a_4249_6147# a_4355_6147# VPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X306 n_d[4].t5 a_5547_7119# VGND.t479 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X307 VGND.t496 _00_ net13 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X308 a_2975_6147# net2 VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X309 VPWR.t364 net1 a_3755_5639# VPWR.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X310 net8 a_4903_6575# VGND.t473 VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X311 VGND.t5 a_4779_7379# n_d[3].t6 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X312 VPWR.t153 VGND.t542 VPWR.t152 VPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X313 net7 a_4745_5533# a_5008_5487# VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X314 n_d[7].t4 a_6099_7119# VGND.t288 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X315 a_5137_2388# in[1].t1 VGND.t251 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X316 a_2387_5461# net16 VPWR.t354 VPWR.t353 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X317 VPWR.t306 _07_ a_4903_6575# VPWR.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X318 VGND.t424 a_2387_5461# y_d[4].t6 VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X319 a_7437_2388# in[2].t0 VPWR.t41 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X320 VGND.t116 VPWR.t524 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X321 VGND.t36 net3 a_4443_3855# VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X322 a_3237_5309# _00_ a_3155_5056# VGND.t494 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X323 a_2667_5175# _00_ VGND.t493 VGND.t492 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X324 VGND.t119 VPWR.t525 VGND.t118 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X325 a_3701_6147# a_3513_6147# a_3619_6147# VPWR.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X326 VPWR.t150 VGND.t543 VPWR.t149 VPWR.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X327 VPWR.t356 a_3019_7338# net18 VPWR.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X328 n_d[2].t0 a_3307_7379# VPWR.t65 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X329 VPWR.t7 a_4779_7379# n_d[3].t3 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X330 VGND.t328 VPWR.t526 VGND.t327 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X331 y_d[4].t5 a_2387_5461# VGND.t422 VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X332 VPWR.t63 _08_ a_3615_4943# VPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X333 VGND.t428 a_3111_5639# _09_ VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X334 VGND.t216 a_3491_6549# y_d[5].t6 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X335 a_3220_4215# net1 a_3148_4215# VGND.t371 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X336 VPWR.t406 a_2387_4373# y_d[3].t1 VPWR.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X337 VPWR.t147 VGND.t544 VPWR.t146 VPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X338 a_3111_5639# a_3384_5467# a_3342_5493# VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X339 VPWR.t475 _00_ a_4745_5533# VPWR.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X340 a_4779_7379# net7 VPWR.t73 VPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X341 VPWR.t144 VGND.t545 VPWR.t143 VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X342 _00_ a_4443_3855# VGND.t284 VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X343 VGND.t337 a_7111_6575# n_d[6].t6 VGND.t336 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X344 VGND.t477 a_5547_7119# n_d[4].t4 VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X345 VGND.t276 a_3219_3463# net13 VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X346 VGND.t331 VPWR.t527 VGND.t330 VGND.t329 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X347 n_d[3].t5 a_4779_7379# VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X348 a_2387_7379# net18 VPWR.t288 VPWR.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X349 VGND.t322 VPWR.t528 VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X350 net10 a_5297_6147# VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X351 VGND.t269 _07_ a_4903_6575# VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X352 a_7437_2388# in[2].t1 VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X353 a_3155_5056# _01_.t18 VPWR.t448 VPWR.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X354 VPWR.t141 VGND.t546 VPWR.t140 VPWR.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X355 y_d[2].t7 a_2387_3027# VGND.t449 VGND.t448 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X356 VPWR.t138 VGND.t547 VPWR.t137 VPWR.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X357 a_4924_5487# _02_ VGND.t389 VGND.t388 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X358 VGND.t370 net1 a_4355_6147# VGND.t369 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X359 VGND.t325 VPWR.t529 VGND.t324 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X360 VGND.t364 net9 a_6651_7119# VGND.t363 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X361 VGND.t135 _08_ a_3615_4943# VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X362 n_d[3].t2 a_4779_7379# VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X363 VGND.t420 a_2387_5461# y_d[4].t4 VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X364 VPWR.t388 _02_ net10 VPWR.t387 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X365 VGND.t491 _00_ net14 VGND.t490 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X366 VGND.t76 VPWR.t530 VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X367 VPWR.t136 VGND.t548 VPWR.t135 VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X368 y_d[5].t5 a_3491_6549# VGND.t214 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X369 VPWR.t133 VGND.t549 VPWR.t132 VPWR.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X370 y_d[3].t0 a_2387_4373# VPWR.t404 VPWR.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X371 y_d[0].t2 a_2879_2223# VPWR.t274 VPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X372 VPWR.t130 VGND.t550 VPWR.t129 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X373 a_5476_6351# _00_ VGND.t489 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X374 VGND.t79 VPWR.t531 VGND.t78 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X375 n_d[6].t5 a_7111_6575# VGND.t335 VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X376 y_d[1].t7 a_2387_2197# VGND.t247 VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X377 VGND.t23 net2 a_3220_4215# VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X378 VGND.t185 VPWR.t532 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X379 VPWR.t127 VGND.t551 VPWR.t126 VPWR.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X380 VGND.t457 _01_.t19 a_3384_5467# VGND.t456 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X381 VPWR.t124 VGND.t552 VPWR.t123 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X382 y_d[0].t6 a_2879_2223# VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X383 VGND.t487 _00_ net12 VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X384 VGND.t21 net2 a_4167_3311# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X385 net16 _02_ VGND.t387 VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X386 a_3773_6147# net1 a_3701_6147# VPWR.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X387 n_d[5].t2 a_6651_7119# VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X388 y_d[6].t6 a_2387_7379# VGND.t300 VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X389 VGND.t188 VPWR.t533 VGND.t187 VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X390 VPWR.t375 net10 a_7111_6575# VPWR.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X391 VGND.t447 a_2387_3027# y_d[2].t6 VGND.t446 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X392 VGND.t110 VPWR.t534 VGND.t109 VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X393 a_2387_3027# net14 VPWR.t377 VPWR.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X394 a_2961_3855# _00_ VGND.t485 VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X395 VGND.t113 VPWR.t535 VGND.t112 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X396 a_5437_6575# _01_.t20 a_5353_6575# VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X397 VPWR.t121 VGND.t553 VPWR.t120 VPWR.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X398 net9 a_5849_6147# VPWR.t381 VPWR.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X399 VGND.t254 VPWR.t536 VGND.t253 VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X400 a_3859_7379# net5 VGND.t408 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X401 y_d[2].t5 a_2387_3027# VGND.t445 VGND.t444 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X402 VPWR.t272 a_2879_2223# y_d[0].t1 VPWR.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X403 VPWR.t47 a_3571_4074# net15 VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X404 VPWR.t386 _02_ a_5849_6147# VPWR.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X405 n_d[3].t1 a_4779_7379# VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X406 VGND.t256 VPWR.t537 VGND.t255 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X407 VGND.t453 a_2376_6263# _03_ VGND.t452 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X408 VPWR.t118 VGND.t554 VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X409 y_d[7].t6 a_2387_6549# VGND.t467 VGND.t466 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X410 VGND.t245 a_2387_2197# y_d[1].t6 VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X411 y_d[5].t4 a_3491_6549# VGND.t212 VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X412 VGND.t316 VPWR.t538 VGND.t315 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X413 VGND.t319 VPWR.t539 VGND.t318 VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X414 VGND.t173 VPWR.t540 VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X415 VPWR.t115 VGND.t555 VPWR.t114 VPWR.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X416 VPWR.t418 a_2387_5461# y_d[4].t2 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X417 VGND.t176 VPWR.t541 VGND.t175 VGND.t174 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X418 VGND.t1 a_4779_7379# n_d[3].t4 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X419 VPWR.t300 _01_.t21 net9 VPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X420 n_d[6].t4 a_7111_6575# VGND.t333 VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X421 y_d[1].t5 a_2387_2197# VGND.t243 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X422 VGND.t223 a_2879_2223# y_d[0].t5 VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X423 VPWR.t49 a_4167_3311# _02_ VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X424 a_4307_6740# _03_ VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X425 y_d[4].t1 a_2387_5461# VPWR.t416 VPWR.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X426 a_3111_5639# a_3384_5467# VPWR.t268 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X427 VPWR.t89 a_6651_7119# n_d[5].t1 VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X428 a_2387_4373# net15 VGND.t182 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X429 a_2376_6263# net3 VGND.t34 VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X430 VPWR.t262 a_3491_6549# y_d[5].t1 VPWR.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X431 VPWR.t473 _00_ a_3155_5056# VPWR.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X432 _07_ a_4355_6147# VPWR.t331 VPWR.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X433 VGND.t298 a_2387_7379# y_d[6].t5 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X434 a_2961_2767# _02_ net12 VPWR.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X435 VGND.t231 a_2939_6549# n_d[0].t4 VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X436 VPWR.t112 VGND.t556 VPWR.t111 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X437 VPWR.t77 net12 a_2879_2223# VPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X438 VPWR.t1 a_4779_7379# n_d[3].t0 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X439 VPWR.t109 VGND.t557 VPWR.t108 VPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X440 y_d[6].t4 a_2387_7379# VGND.t296 VGND.t295 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X441 VGND.t443 a_2387_3027# y_d[2].t4 VGND.t442 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X442 y_d[0].t0 a_2879_2223# VPWR.t270 VPWR.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X443 a_2387_6549# net19 VPWR.t361 VPWR.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X444 VGND.t465 a_2387_6549# y_d[7].t5 VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X445 VPWR.t325 a_2387_7379# y_d[6].t1 VPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X446 VGND.t279 VPWR.t542 VGND.t278 VGND.t277 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X447 VGND.t282 VPWR.t543 VGND.t281 VGND.t280 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X448 net9 _00_ VPWR.t471 VPWR.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X449 a_2511_6147# net3 VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X450 a_3619_6147# net1 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X451 VGND.t103 VPWR.t544 VGND.t102 VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X452 y_d[7].t4 a_2387_6549# VGND.t463 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X453 n_d[0].t0 a_2939_6549# VPWR.t280 VPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X454 VPWR.t106 VGND.t558 VPWR.t105 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X455 a_3219_3463# _01_.t22 VGND.t180 VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X456 a_3219_3463# _01_.t23 VPWR.t81 VPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X457 VGND.t106 VPWR.t545 VGND.t105 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X458 y_d[6].t0 a_2387_7379# VPWR.t323 VPWR.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X459 VGND.t241 a_2387_2197# y_d[1].t4 VGND.t240 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X460 y_d[0].t4 a_2879_2223# VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X461 VGND.t155 VPWR.t546 VGND.t154 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X462 _04_ a_2975_6147# VGND.t431 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X463 VPWR.t103 VGND.t559 VPWR.t102 VPWR.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X464 a_4307_6740# _03_ VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X465 VPWR.t414 a_2387_5461# y_d[4].t0 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X466 VGND.t11 a_2667_5175# net16 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X467 VGND.t158 VPWR.t547 VGND.t157 VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X468 n_d[5].t0 a_6651_7119# VPWR.t87 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X469 VPWR.t100 VGND.t560 VPWR.t99 VPWR.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X470 net11 _02_ VPWR.t383 VPWR.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X471 y_d[5].t0 a_3491_6549# VPWR.t260 VPWR.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R0 VGND.n1191 VGND 4653.9
R1 VGND VGND.n839 4242.17
R2 VGND.n836 VGND 4140.08
R3 VGND.t165 VGND 4121.84
R4 VGND.t174 VGND 4121.84
R5 VGND.n837 VGND.n836 3873.14
R6 VGND.n838 VGND.n837 3873.14
R7 VGND.n839 VGND.n838 3873.14
R8 VGND VGND.t329 3632.95
R9 VGND VGND.t189 3632.95
R10 VGND.n1194 VGND 3595.55
R11 VGND.t74 VGND.t86 3101.92
R12 VGND.t129 VGND.t252 3101.92
R13 VGND.t317 VGND.n383 2714.18
R14 VGND.t12 VGND.t83 2714.18
R15 VGND.t48 VGND.t171 2714.18
R16 VGND.t257 VGND 2570.88
R17 VGND VGND.t120 2562.45
R18 VGND VGND.t126 2452.87
R19 VGND.n1194 VGND.n1193 2410.47
R20 VGND.n1193 VGND.n1192 2410.47
R21 VGND.n1192 VGND.n1191 2410.47
R22 VGND.t120 VGND.t186 2326.44
R23 VGND.t89 VGND.t317 2326.44
R24 VGND.t150 VGND.t257 2326.44
R25 VGND VGND.t89 2081.99
R26 VGND VGND.t150 2081.99
R27 VGND VGND.t114 2081.99
R28 VGND.t338 VGND.t15 2022.99
R29 VGND.t452 VGND.t262 1989.27
R30 VGND.t86 VGND 1795.4
R31 VGND.t252 VGND 1795.4
R32 VGND VGND.n547 1677.39
R33 VGND.t399 VGND.t239 1576.25
R34 VGND.t429 VGND.t484 1576.25
R35 VGND.t65 VGND.t153 1567.82
R36 VGND.n384 VGND.t117 1550.96
R37 VGND.t280 VGND.t77 1550.96
R38 VGND VGND.t385 1458.24
R39 VGND.t73 VGND 1458.24
R40 VGND VGND.t179 1432.95
R41 VGND VGND.t111 1407.66
R42 VGND VGND.t168 1407.66
R43 VGND VGND.t95 1407.66
R44 VGND VGND.t326 1306.51
R45 VGND VGND.t12 1306.51
R46 VGND.t171 VGND 1306.51
R47 VGND VGND.t74 1306.51
R48 VGND VGND.t129 1306.51
R49 VGND.t427 VGND.t492 1205.36
R50 VGND.n1318 VGND.n24 1198.25
R51 VGND.n183 VGND.n182 1198.25
R52 VGND.n549 VGND.n548 1198.25
R53 VGND.n841 VGND.n840 1198.25
R54 VGND.n1190 VGND.n1189 1198.25
R55 VGND.n835 VGND.n834 1198.25
R56 VGND.n1089 VGND.n993 1194.5
R57 VGND.n1196 VGND.n1195 1194.5
R58 VGND.n383 VGND.n382 1194.5
R59 VGND.n697 VGND.n384 1194.5
R60 VGND.n547 VGND.n546 1194.5
R61 VGND.n992 VGND.n991 1194.5
R62 VGND VGND.t156 1048.99
R63 VGND VGND.t472 1028.35
R64 VGND VGND.t69 1028.35
R65 VGND VGND.t61 1028.35
R66 VGND.t114 VGND 1019.92
R67 VGND VGND.t280 1011.49
R68 VGND.t37 VGND.t207 977.779
R69 VGND.t474 VGND.t22 977.779
R70 VGND.t156 VGND 944.277
R71 VGND VGND.n992 927.203
R72 VGND.n993 VGND 927.203
R73 VGND.t262 VGND 918.774
R74 VGND.t111 VGND 918.774
R75 VGND.t168 VGND 918.774
R76 VGND.t95 VGND 918.774
R77 VGND.t385 VGND.t270 901.917
R78 VGND.t47 VGND.t396 901.917
R79 VGND VGND.t73 868.199
R80 VGND.n836 VGND 851.341
R81 VGND.n837 VGND 851.341
R82 VGND.n838 VGND 851.341
R83 VGND.n839 VGND 851.341
R84 VGND.t232 VGND.t373 842.913
R85 VGND.t405 VGND.t460 834.484
R86 VGND.t500 VGND.t388 817.625
R87 VGND.t492 VGND.t313 817.625
R88 VGND.t181 VGND.t413 817.625
R89 VGND.t179 VGND.t495 817.625
R90 VGND.t498 VGND 809.196
R91 VGND.t430 VGND.t234 800.766
R92 VGND.t18 VGND.t219 800.766
R93 VGND.t67 VGND.t20 800.766
R94 VGND.t63 VGND.t375 800.766
R95 VGND.t438 VGND.t39 775.48
R96 VGND.t456 VGND.t18 775.48
R97 VGND.t329 VGND.t165 775.48
R98 VGND.t189 VGND.t174 775.48
R99 VGND.t403 VGND 767.051
R100 VGND VGND.t500 767.051
R101 VGND.n840 VGND.t162 747.476
R102 VGND.t228 VGND.t432 741.763
R103 VGND.t472 VGND.t268 741.763
R104 VGND.t8 VGND.t438 741.763
R105 VGND.t99 VGND.t134 741.763
R106 VGND.t458 VGND.t65 741.763
R107 VGND.t336 VGND.t334 724.904
R108 VGND.t213 VGND.t215 724.904
R109 VGND.t215 VGND.t211 724.904
R110 VGND.t230 VGND.t232 724.904
R111 VGND.t468 VGND.t462 724.904
R112 VGND.t425 VGND.t419 724.904
R113 VGND.t415 VGND.t409 724.904
R114 VGND.t409 VGND.t411 724.904
R115 VGND.t448 VGND.t442 724.904
R116 VGND.t342 VGND 720.394
R117 VGND.t270 VGND.t498 708.047
R118 VGND.t41 VGND.t367 708.047
R119 VGND.t43 VGND.t24 708.047
R120 VGND.t24 VGND.t434 708.047
R121 VGND.t388 VGND.t249 708.047
R122 VGND.t413 VGND.t123 708.047
R123 VGND.t61 VGND.t63 708.047
R124 VGND.t495 VGND.t397 708.047
R125 VGND.t397 VGND.t275 708.047
R126 VGND.t486 VGND.t271 708.047
R127 VGND.t104 VGND.t338 691.188
R128 VGND.t22 VGND.t371 682.76
R129 VGND.t464 VGND.t377 674.331
R130 VGND.t217 VGND.t450 657.471
R131 VGND.t466 VGND.t33 657.471
R132 VGND.t372 VGND 657.471
R133 VGND VGND.t386 649.043
R134 VGND VGND.t311 640.614
R135 VGND.t15 VGND 632.184
R136 VGND.t126 VGND 632.184
R137 VGND.n383 VGND 632.184
R138 VGND.n384 VGND 632.184
R139 VGND.t83 VGND 632.184
R140 VGND VGND.t48 632.184
R141 VGND.n993 VGND 632.184
R142 VGND.t421 VGND 615.327
R143 VGND.t411 VGND 615.327
R144 VGND.t444 VGND 615.327
R145 VGND.t162 VGND 612.064
R146 VGND VGND.t342 612.064
R147 VGND.t239 VGND.t372 606.898
R148 VGND.t371 VGND.t429 606.898
R149 VGND.t283 VGND 590.038
R150 VGND VGND.n1194 564.751
R151 VGND.n1193 VGND 564.751
R152 VGND.n1192 VGND 564.751
R153 VGND.n1191 VGND 564.751
R154 VGND.t379 VGND 556.322
R155 VGND.t35 VGND 556.322
R156 VGND.t20 VGND 556.322
R157 VGND VGND.t336 547.894
R158 VGND.t39 VGND 547.894
R159 VGND.t28 VGND 547.894
R160 VGND.t373 VGND 547.894
R161 VGND.t134 VGND 547.894
R162 VGND.t494 VGND 547.894
R163 VGND.t392 VGND 539.465
R164 VGND.t484 VGND 539.465
R165 VGND.t58 VGND.t277 535.653
R166 VGND.t186 VGND 531.034
R167 VGND.t303 VGND 531.034
R168 VGND.t159 VGND 531.034
R169 VGND.t77 VGND 531.034
R170 VGND.t306 VGND 531.034
R171 VGND.t205 VGND 522.606
R172 VGND.t10 VGND.t423 522.606
R173 VGND.t436 VGND.t446 522.606
R174 VGND.t30 VGND 514.177
R175 VGND.t69 VGND 514.177
R176 VGND.t132 VGND.t80 501.93
R177 VGND.t365 VGND 497.318
R178 VGND.t248 VGND.t273 488.889
R179 VGND.t460 VGND 488.889
R180 VGND.t497 VGND.t488 480.461
R181 VGND.n1195 VGND.t369 472.031
R182 VGND.t390 VGND.t490 472.031
R183 VGND.t423 VGND 463.603
R184 VGND.t446 VGND 463.603
R185 VGND.n182 VGND.t332 455.173
R186 VGND.t432 VGND.t47 455.173
R187 VGND.t369 VGND 455.173
R188 VGND.t183 VGND.t242 433.32
R189 VGND.t419 VGND.t320 421.457
R190 VGND.t442 VGND.t101 421.457
R191 VGND.t98 VGND.t45 404.599
R192 VGND.t192 VGND.t295 399.245
R193 VGND.t117 VGND.t159 387.74
R194 VGND.n547 VGND.t55 387.74
R195 VGND.n992 VGND.t265 387.74
R196 VGND.n548 VGND.t285 370.882
R197 VGND VGND.t92 366.517
R198 VGND.n182 VGND.t379 362.452
R199 VGND VGND.t486 362.452
R200 VGND.t271 VGND.t401 362.452
R201 VGND VGND.n1190 359.295
R202 VGND.n1195 VGND.t309 345.594
R203 VGND.t401 VGND.t390 345.594
R204 VGND.n548 VGND.t283 337.166
R205 VGND.t488 VGND.t248 328.736
R206 VGND.t394 VGND.t32 328.736
R207 VGND VGND.t309 303.449
R208 VGND.t320 VGND.t421 303.449
R209 VGND.t101 VGND.t444 303.449
R210 VGND.t357 VGND.t10 295.019
R211 VGND.t381 VGND.t436 295.019
R212 VGND VGND.t26 286.591
R213 VGND VGND.t417 285.269
R214 VGND.t80 VGND 279.853
R215 VGND.n1057 VGND.t487 278.589
R216 VGND.t219 VGND.t394 278.161
R217 VGND.t32 VGND.t98 278.161
R218 VGND VGND.t323 277.808
R219 VGND.n957 VGND.t559 276.101
R220 VGND.n209 VGND.t393 274.812
R221 VGND VGND.t353 274.481
R222 VGND VGND.t142 274.481
R223 VGND VGND.t454 269.733
R224 VGND VGND.t440 269.733
R225 VGND VGND.t365 269.733
R226 VGND VGND.t357 269.733
R227 VGND VGND.t181 269.733
R228 VGND VGND.t381 269.733
R229 VGND.n1090 VGND.t522 265.298
R230 VGND VGND.t359 262.837
R231 VGND.n793 VGND.t523 262.784
R232 VGND.n794 VGND.t529 262.784
R233 VGND.n1226 VGND.t507 262.784
R234 VGND.n1228 VGND.t514 262.784
R235 VGND.n636 VGND.t550 262.784
R236 VGND.n638 VGND.t552 262.784
R237 VGND.n342 VGND.t506 262.784
R238 VGND.n358 VGND.t510 262.784
R239 VGND.n576 VGND.t535 262.784
R240 VGND.n577 VGND.t537 262.784
R241 VGND.n416 VGND.t548 262.784
R242 VGND.n417 VGND.t551 262.784
R243 VGND.n146 VGND.t533 262.784
R244 VGND.n147 VGND.t536 262.784
R245 VGND.n1031 VGND.t518 262.784
R246 VGND.n1033 VGND.t519 262.784
R247 VGND.n936 VGND.t541 262.719
R248 VGND.n141 VGND.t504 262.719
R249 VGND.n195 VGND.t505 262.719
R250 VGND.n388 VGND.t540 262.719
R251 VGND.n371 VGND.t508 262.719
R252 VGND.n742 VGND.t531 262.719
R253 VGND.n317 VGND.t528 262.719
R254 VGND.n318 VGND.t539 262.719
R255 VGND.n496 VGND.t520 262.719
R256 VGND.n470 VGND.t553 262.719
R257 VGND.n519 VGND.t556 262.719
R258 VGND.n521 VGND.t534 262.719
R259 VGND.n600 VGND.t516 262.719
R260 VGND.n123 VGND.t512 262.719
R261 VGND.n1012 VGND.t543 262.719
R262 VGND VGND.t228 261.303
R263 VGND VGND.t205 261.303
R264 VGND.t326 VGND 261.303
R265 VGND VGND.t425 261.303
R266 VGND.t285 VGND 261.303
R267 VGND VGND.t458 261.303
R268 VGND VGND.t448 261.303
R269 VGND VGND.t361 261.173
R270 VGND.n1222 VGND.t374 259.51
R271 VGND.n1277 VGND.t40 259.51
R272 VGND.n675 VGND.t457 259.51
R273 VGND.n1357 VGND.t513 259.082
R274 VGND.n265 VGND.t549 259.082
R275 VGND.n643 VGND.t544 259.082
R276 VGND.n692 VGND.t554 259.082
R277 VGND.n160 VGND.t517 259.082
R278 VGND.n87 VGND.t557 259.082
R279 VGND.n1038 VGND.t511 259.082
R280 VGND.n820 VGND.t526 259.082
R281 VGND.t277 VGND 257.846
R282 VGND.n1218 VGND.t29 255.326
R283 VGND.n689 VGND.t400 255.326
R284 VGND.n592 VGND.t485 255.326
R285 VGND VGND.t30 252.875
R286 VGND VGND.t399 252.875
R287 VGND VGND.t456 252.875
R288 VGND.n835 VGND.t197 246.201
R289 VGND.t6 VGND.n24 246.201
R290 VGND.t55 VGND 244.445
R291 VGND VGND.t265 244.445
R292 VGND.n1353 VGND.t296 243.286
R293 VGND.n1348 VGND.t143 243.286
R294 VGND.n16 VGND.t354 243.286
R295 VGND.n23 VGND.t7 243.286
R296 VGND.n280 VGND.t481 243.286
R297 VGND.n249 VGND.t294 243.286
R298 VGND.n163 VGND.t198 243.286
R299 VGND.n1230 VGND.t463 243.286
R300 VGND.n1243 VGND.t233 243.286
R301 VGND.n108 VGND.t227 243.286
R302 VGND.n83 VGND.t243 243.286
R303 VGND.t226 VGND 240.131
R304 VGND.n179 VGND.t339 239.4
R305 VGND.n1206 VGND.t212 239.4
R306 VGND.n642 VGND.t422 239.4
R307 VGND.n580 VGND.t412 239.4
R308 VGND.n1037 VGND.t445 239.4
R309 VGND.n413 VGND.t286 238.558
R310 VGND.n1000 VGND.t62 235.607
R311 VGND.n1084 VGND.t70 235.607
R312 VGND.t396 VGND.t497 227.587
R313 VGND VGND.t427 227.587
R314 VGND.n362 VGND.t542 224.094
R315 VGND.n513 VGND.t331 223.662
R316 VGND.n448 VGND.t166 223.438
R317 VGND.n466 VGND.t175 223.438
R318 VGND.t209 VGND 222.077
R319 VGND.n484 VGND.t191 220.16
R320 VGND.t273 VGND.t392 219.157
R321 VGND VGND.t405 219.157
R322 VGND.n786 VGND.t560 218.308
R323 VGND.n44 VGND.t532 218.308
R324 VGND.n440 VGND.t525 218.308
R325 VGND.n1119 VGND.t545 218.308
R326 VGND.n911 VGND.t509 218.308
R327 VGND.n829 VGND.t558 218.308
R328 VGND.n338 VGND.t318 217.977
R329 VGND.n408 VGND.t154 217.977
R330 VGND VGND.t293 217.922
R331 VGND VGND.t480 217.922
R332 VGND.n184 VGND.t121 216.933
R333 VGND.n985 VGND.t115 215.992
R334 VGND.n362 VGND.t328 214.488
R335 VGND.n1356 VGND.t194 214.456
R336 VGND.n1359 VGND.t193 214.456
R337 VGND.n821 VGND.t60 214.456
R338 VGND.n819 VGND.t59 214.456
R339 VGND.n165 VGND.t279 214.456
R340 VGND.n827 VGND.t278 214.456
R341 VGND.n264 VGND.t325 214.456
R342 VGND.n267 VGND.t324 214.456
R343 VGND.n917 VGND.t267 214.456
R344 VGND.n919 VGND.t87 214.456
R345 VGND.n979 VGND.t116 214.456
R346 VGND.n937 VGND.t88 214.456
R347 VGND.n928 VGND.t75 214.456
R348 VGND.n938 VGND.t253 214.456
R349 VGND.n951 VGND.t76 214.456
R350 VGND.n143 VGND.t254 214.456
R351 VGND.n942 VGND.t130 214.456
R352 VGND.n1083 VGND.t131 214.456
R353 VGND.n1059 VGND.t308 214.456
R354 VGND.n997 VGND.t307 214.456
R355 VGND.n785 VGND.t106 214.456
R356 VGND.n177 VGND.t105 214.456
R357 VGND.n793 VGND.t341 214.456
R358 VGND.n793 VGND.t340 214.456
R359 VGND.n794 VGND.t17 214.456
R360 VGND.n794 VGND.t16 214.456
R361 VGND.n48 VGND.t305 214.456
R362 VGND.n43 VGND.t304 214.456
R363 VGND.n1226 VGND.t316 214.456
R364 VGND.n1226 VGND.t315 214.456
R365 VGND.n1228 VGND.t264 214.456
R366 VGND.n1228 VGND.t263 214.456
R367 VGND.n198 VGND.t188 214.456
R368 VGND.n765 VGND.t122 214.456
R369 VGND.n775 VGND.t187 214.456
R370 VGND.n319 VGND.t259 214.456
R371 VGND.n313 VGND.t151 214.456
R372 VGND.n329 VGND.t152 214.456
R373 VGND.n336 VGND.t160 214.456
R374 VGND.n691 VGND.t119 214.456
R375 VGND.n387 VGND.t118 214.456
R376 VGND.n390 VGND.t161 214.456
R377 VGND.n641 VGND.t322 214.456
R378 VGND.n634 VGND.t321 214.456
R379 VGND.n636 VGND.t149 214.456
R380 VGND.n636 VGND.t148 214.456
R381 VGND.n638 VGND.t113 214.456
R382 VGND.n638 VGND.t112 214.456
R383 VGND.n312 VGND.t258 214.456
R384 VGND.n728 VGND.t91 214.456
R385 VGND.n741 VGND.t319 214.456
R386 VGND.n368 VGND.t90 214.456
R387 VGND.n361 VGND.t327 214.456
R388 VGND.n342 VGND.t256 214.456
R389 VGND.n342 VGND.t255 214.456
R390 VGND.n358 VGND.t128 214.456
R391 VGND.n358 VGND.t127 214.456
R392 VGND.n576 VGND.t261 214.456
R393 VGND.n576 VGND.t260 214.456
R394 VGND.n577 VGND.t170 214.456
R395 VGND.n577 VGND.t169 214.456
R396 VGND.n573 VGND.t124 214.456
R397 VGND.n584 VGND.t125 214.456
R398 VGND.n594 VGND.t155 214.456
R399 VGND.n562 VGND.t79 214.456
R400 VGND.n409 VGND.t282 214.456
R401 VGND.n559 VGND.t78 214.456
R402 VGND.n553 VGND.t281 214.456
R403 VGND.n437 VGND.t56 214.456
R404 VGND.n439 VGND.t14 214.456
R405 VGND.n437 VGND.t13 214.456
R406 VGND.n416 VGND.t85 214.456
R407 VGND.n416 VGND.t84 214.456
R408 VGND.n417 VGND.t110 214.456
R409 VGND.n417 VGND.t109 214.456
R410 VGND.n447 VGND.t57 214.456
R411 VGND.n536 VGND.t330 214.456
R412 VGND.n465 VGND.t167 214.456
R413 VGND.n508 VGND.t190 214.456
R414 VGND.n483 VGND.t176 214.456
R415 VGND.n86 VGND.t185 214.456
R416 VGND.n89 VGND.t184 214.456
R417 VGND.n57 VGND.t344 214.456
R418 VGND.n1183 VGND.t343 214.456
R419 VGND.n1118 VGND.t82 214.456
R420 VGND.n129 VGND.t81 214.456
R421 VGND.n125 VGND.t158 214.456
R422 VGND.n120 VGND.t157 214.456
R423 VGND.n847 VGND.t164 214.456
R424 VGND.n868 VGND.t163 214.456
R425 VGND.n880 VGND.t94 214.456
R426 VGND.n159 VGND.t93 214.456
R427 VGND.n908 VGND.t266 214.456
R428 VGND.n910 VGND.t173 214.456
R429 VGND.n908 VGND.t172 214.456
R430 VGND.n146 VGND.t52 214.456
R431 VGND.n146 VGND.t51 214.456
R432 VGND.n147 VGND.t50 214.456
R433 VGND.n147 VGND.t49 214.456
R434 VGND.n1036 VGND.t103 214.456
R435 VGND.n1029 VGND.t102 214.456
R436 VGND.n1031 VGND.t97 214.456
R437 VGND.n1031 VGND.t96 214.456
R438 VGND.n1033 VGND.t346 214.456
R439 VGND.n1033 VGND.t345 214.456
R440 VGND VGND.t35 210.728
R441 VGND.t275 VGND 210.728
R442 VGND.n396 VGND.n395 208.553
R443 VGND.n1366 VGND.n1365 205.078
R444 VGND.n2 VGND.n1 205.078
R445 VGND.n1329 VGND.n18 205.078
R446 VGND.n1313 VGND.n27 205.078
R447 VGND.n276 VGND.n275 205.078
R448 VGND.n295 VGND.n294 205.078
R449 VGND.n243 VGND.n239 205.078
R450 VGND.n1224 VGND.n1223 205.078
R451 VGND.n1265 VGND.n1264 205.078
R452 VGND.n106 VGND.n75 205.078
R453 VGND.n95 VGND.n82 205.078
R454 VGND.n1247 VGND.n1245 204.109
R455 VGND.n1351 VGND.n1350 203.619
R456 VGND.n1335 VGND.n15 203.619
R457 VGND.n20 VGND.n19 203.619
R458 VGND.n29 VGND.n28 203.619
R459 VGND.n273 VGND.n272 203.619
R460 VGND.n283 VGND.n282 203.619
R461 VGND.n237 VGND.n236 203.619
R462 VGND.n1239 VGND.n1238 203.619
R463 VGND.n1204 VGND.n1203 203.619
R464 VGND.n412 VGND.n411 203.619
R465 VGND.n78 VGND.n77 203.619
R466 VGND.n80 VGND.n79 203.619
R467 VGND.n183 VGND.n181 203.415
R468 VGND.n662 VGND.n627 203.22
R469 VGND.n679 VGND.n393 203.22
R470 VGND.n1252 VGND.n1220 202.564
R471 VGND.n204 VGND.n203 202.349
R472 VGND.t45 VGND.t494 202.299
R473 VGND.n787 VGND.n180 200.812
R474 VGND.n648 VGND.n633 200.812
R475 VGND.n580 VGND.n579 200.812
R476 VGND.n1043 VGND.n1028 200.812
R477 VGND.n767 VGND.n766 200.692
R478 VGND.n1174 VGND.n56 200.692
R479 VGND.n859 VGND.n846 200.692
R480 VGND.n1237 VGND.n1236 200.516
R481 VGND.n1247 VGND.n1246 200.516
R482 VGND.n1267 VGND.n1266 200.516
R483 VGND.n1283 VGND.n1282 200.516
R484 VGND.n569 VGND.n568 199.917
R485 VGND.n1377 VGND.n1376 199.739
R486 VGND.n22 VGND.n21 199.739
R487 VGND.n1202 VGND.n1201 199.739
R488 VGND.n1200 VGND.n1199 199.739
R489 VGND.n200 VGND.n199 199.739
R490 VGND.n392 VGND.n391 199.739
R491 VGND.n162 VGND.n161 199.739
R492 VGND.n127 VGND.n126 199.739
R493 VGND.n59 VGND.n58 199.739
R494 VGND.n1073 VGND.n1001 199.662
R495 VGND.n1081 VGND.n996 199.662
R496 VGND.n650 VGND.n632 199.662
R497 VGND.n587 VGND.n575 199.662
R498 VGND.n1045 VGND.n1027 199.662
R499 VGND.n197 VGND.n196 199.052
R500 VGND.n337 VGND.n328 199.052
R501 VGND.n1252 VGND.n1251 198.654
R502 VGND.n1272 VGND.n1271 198.654
R503 VGND.n1232 VGND.n1231 198.475
R504 VGND.n630 VGND.n629 196.831
R505 VGND.n1025 VGND.n1024 196.831
R506 VGND.n1052 VGND.n1022 196.831
R507 VGND.n1060 VGND.n1019 196.831
R508 VGND VGND.t183 196.799
R509 VGND.n1297 VGND.n42 196.442
R510 VGND.n567 VGND.n406 196.442
R511 VGND.n1198 VGND.n1197 195.752
R512 VGND VGND.t502 193.87
R513 VGND VGND.t67 193.87
R514 VGND.n190 VGND.n188 190.399
R515 VGND.n1176 VGND.n1175 190.399
R516 VGND.n861 VGND.n860 190.399
R517 VGND.t323 VGND 181.323
R518 VGND VGND.n24 181.323
R519 VGND VGND.t192 181.323
R520 VGND.t332 VGND 177.012
R521 VGND.t146 VGND.t224 175.133
R522 VGND.t244 VGND.t470 175.133
R523 VGND.t203 VGND.t363 161.362
R524 VGND.t291 VGND.t107 161.362
R525 VGND.t478 VGND.t177 161.362
R526 VGND.t144 VGND.t0 161.362
R527 VGND.t349 VGND.t407 161.362
R528 VGND.t138 VGND.t355 161.362
R529 VGND.t297 VGND.t237 161.362
R530 VGND.t417 VGND.t53 158.885
R531 VGND.t250 VGND.t132 158.885
R532 VGND.t71 VGND.t209 158.885
R533 VGND.t220 VGND.t226 155.274
R534 VGND.t222 VGND.t220 155.274
R535 VGND.t224 VGND.t222 155.274
R536 VGND.t246 VGND.t244 155.274
R537 VGND.t240 VGND.t246 155.274
R538 VGND.t242 VGND.t240 155.274
R539 VGND.n768 VGND.n767 152
R540 VGND.n859 VGND.n858 152
R541 VGND.n1174 VGND.n1173 152
R542 VGND.t361 VGND.t383 146.389
R543 VGND.t359 VGND.t195 146.389
R544 VGND.t386 VGND 143.296
R545 VGND.t311 VGND 143.296
R546 VGND.t197 VGND.t199 143.062
R547 VGND.t199 VGND.t201 143.062
R548 VGND.t201 VGND.t203 143.062
R549 VGND.t293 VGND.t287 143.062
R550 VGND.t287 VGND.t289 143.062
R551 VGND.t289 VGND.t291 143.062
R552 VGND.t480 VGND.t482 143.062
R553 VGND.t482 VGND.t476 143.062
R554 VGND.t476 VGND.t478 143.062
R555 VGND.t0 VGND.t2 143.062
R556 VGND.t2 VGND.t4 143.062
R557 VGND.t4 VGND.t6 143.062
R558 VGND.t347 VGND.t349 143.062
R559 VGND.t351 VGND.t347 143.062
R560 VGND.t353 VGND.t351 143.062
R561 VGND.t140 VGND.t138 143.062
R562 VGND.t136 VGND.t140 143.062
R563 VGND.t142 VGND.t136 143.062
R564 VGND.t299 VGND.t297 143.062
R565 VGND.t301 VGND.t299 143.062
R566 VGND.t295 VGND.t301 143.062
R567 VGND.t92 VGND 135.412
R568 VGND.n1190 VGND 135.412
R569 VGND.n840 VGND 133.607
R570 VGND VGND.t58 124.764
R571 VGND VGND.n835 124.764
R572 VGND.n584 VGND.t527 121.927
R573 VGND.n409 VGND.t515 119.645
R574 VGND VGND.t146 119.163
R575 VGND.n980 VGND.t555 116.734
R576 VGND VGND.t71 113.746
R577 VGND.n657 VGND.n656 111.15
R578 VGND.n560 VGND.t546 110.102
R579 VGND.t363 VGND 109.793
R580 VGND.t107 VGND 109.793
R581 VGND.t177 VGND 109.793
R582 VGND.n1051 VGND.n1023 107.853
R583 VGND.n1011 VGND.n1010 107.853
R584 VGND.n395 VGND.t395 101.43
R585 VGND.n446 VGND.t538 94.9001
R586 VGND.n916 VGND.t521 94.6788
R587 VGND.n568 VGND.t23 83.899
R588 VGND.n627 VGND.t46 83.8933
R589 VGND.n393 VGND.t38 83.8933
R590 VGND.t502 VGND.t8 67.4335
R591 VGND.t450 VGND.t213 67.4335
R592 VGND.t211 VGND.t28 67.4335
R593 VGND.t33 VGND.t468 67.4335
R594 VGND.t490 VGND 67.4335
R595 VGND.t454 VGND.t41 59.0043
R596 VGND.t313 VGND 59.0043
R597 VGND.n196 VGND.t404 58.5719
R598 VGND.n203 VGND.t274 58.5719
R599 VGND.n328 VGND.t501 58.5719
R600 VGND.n656 VGND.t493 57.875
R601 VGND.n1023 VGND.t402 57.875
R602 VGND.n1010 VGND.t180 57.875
R603 VGND.t470 VGND 57.7765
R604 VGND.n1350 VGND.t298 55.7148
R605 VGND.n15 VGND.t139 55.7148
R606 VGND.n19 VGND.t350 55.7148
R607 VGND.n28 VGND.t1 55.7148
R608 VGND.n272 VGND.t479 55.7148
R609 VGND.n282 VGND.t292 55.7148
R610 VGND.n236 VGND.t204 55.7148
R611 VGND.n181 VGND.t333 55.7148
R612 VGND.n1238 VGND.t465 55.7148
R613 VGND.n1220 VGND.t235 55.7148
R614 VGND.n1203 VGND.t218 55.7148
R615 VGND.n632 VGND.t424 55.7148
R616 VGND.n575 VGND.t414 55.7148
R617 VGND.n77 VGND.t225 55.7148
R618 VGND.n79 VGND.t245 55.7148
R619 VGND.n1027 VGND.t447 55.7148
R620 VGND VGND.t144 53.233
R621 VGND.t407 VGND 53.233
R622 VGND.t355 VGND 53.233
R623 VGND.t237 VGND 53.233
R624 VGND.n1001 VGND.t64 52.8576
R625 VGND.n996 VGND.t68 52.8576
R626 VGND.n1231 VGND.t34 52.8576
R627 VGND.n411 VGND.t284 52.8576
R628 VGND.t53 VGND 52.36
R629 VGND VGND.t250 52.36
R630 VGND.t383 VGND 51.5695
R631 VGND.t195 VGND 51.5695
R632 VGND.n1251 VGND.t44 51.4291
R633 VGND.n1271 VGND.t42 51.4291
R634 VGND.n1197 VGND.t370 51.4291
R635 VGND.t367 VGND.t217 50.5752
R636 VGND.t377 VGND.t466 50.5752
R637 VGND.n447 VGND.n446 41.557
R638 VGND.n1365 VGND.t300 40.0005
R639 VGND.n1365 VGND.t302 40.0005
R640 VGND.n1350 VGND.t238 40.0005
R641 VGND.n1 VGND.t141 40.0005
R642 VGND.n1 VGND.t137 40.0005
R643 VGND.n15 VGND.t356 40.0005
R644 VGND.n18 VGND.t348 40.0005
R645 VGND.n18 VGND.t352 40.0005
R646 VGND.n19 VGND.t408 40.0005
R647 VGND.n27 VGND.t3 40.0005
R648 VGND.n27 VGND.t5 40.0005
R649 VGND.n28 VGND.t145 40.0005
R650 VGND.n272 VGND.t178 40.0005
R651 VGND.n275 VGND.t483 40.0005
R652 VGND.n275 VGND.t477 40.0005
R653 VGND.n282 VGND.t108 40.0005
R654 VGND.n294 VGND.t288 40.0005
R655 VGND.n294 VGND.t290 40.0005
R656 VGND.n236 VGND.t364 40.0005
R657 VGND.n239 VGND.t200 40.0005
R658 VGND.n239 VGND.t202 40.0005
R659 VGND.n1001 VGND.t376 40.0005
R660 VGND.n996 VGND.t21 40.0005
R661 VGND.n180 VGND.t335 40.0005
R662 VGND.n180 VGND.t337 40.0005
R663 VGND.n181 VGND.t380 40.0005
R664 VGND.n1223 VGND.t467 40.0005
R665 VGND.n1223 VGND.t469 40.0005
R666 VGND.n1238 VGND.t366 40.0005
R667 VGND.n1245 VGND.t236 40.0005
R668 VGND.n1245 VGND.t231 40.0005
R669 VGND.n1220 VGND.t441 40.0005
R670 VGND.n1264 VGND.t214 40.0005
R671 VGND.n1264 VGND.t216 40.0005
R672 VGND.n1203 VGND.t455 40.0005
R673 VGND.n633 VGND.t426 40.0005
R674 VGND.n633 VGND.t420 40.0005
R675 VGND.n632 VGND.t358 40.0005
R676 VGND.n579 VGND.t416 40.0005
R677 VGND.n579 VGND.t410 40.0005
R678 VGND.n411 VGND.t36 40.0005
R679 VGND.n575 VGND.t182 40.0005
R680 VGND.n75 VGND.t221 40.0005
R681 VGND.n75 VGND.t223 40.0005
R682 VGND.n77 VGND.t147 40.0005
R683 VGND.n79 VGND.t471 40.0005
R684 VGND.n82 VGND.t247 40.0005
R685 VGND.n82 VGND.t241 40.0005
R686 VGND.n1028 VGND.t449 40.0005
R687 VGND.n1028 VGND.t443 40.0005
R688 VGND.n1027 VGND.t382 40.0005
R689 VGND.n1236 VGND.t27 38.5719
R690 VGND.n1236 VGND.t378 38.5719
R691 VGND.n1246 VGND.t25 38.5719
R692 VGND.n1246 VGND.t435 38.5719
R693 VGND.n1266 VGND.t368 38.5719
R694 VGND.n1266 VGND.t451 38.5719
R695 VGND.n1282 VGND.t31 38.5719
R696 VGND.n1282 VGND.t503 38.5719
R697 VGND.n1372 VGND.n1349 34.6358
R698 VGND.n1372 VGND.n1371 34.6358
R699 VGND.n1324 VGND.n1323 34.6358
R700 VGND.n1288 VGND.n1196 34.6358
R701 VGND.n215 VGND.n214 34.6358
R702 VGND.n214 VGND.n201 34.6358
R703 VGND.n655 VGND.n654 34.6358
R704 VGND.n658 VGND.n626 34.6358
R705 VGND.n664 VGND.n663 34.6358
R706 VGND.n874 VGND.n873 34.6358
R707 VGND.n1188 VGND.n51 34.6358
R708 VGND.n101 VGND.n100 34.6358
R709 VGND.n1050 VGND.n1049 34.6358
R710 VGND.n1053 VGND.n1020 34.6358
R711 VGND.n190 VGND.t530 34.2973
R712 VGND.n1175 VGND.t524 34.2973
R713 VGND.n860 VGND.t547 34.2973
R714 VGND.n650 VGND.n649 34.2593
R715 VGND.n1045 VGND.n1044 34.2593
R716 VGND.t334 VGND.t104 33.717
R717 VGND.t26 VGND.t464 33.717
R718 VGND.t462 VGND.t452 33.717
R719 VGND.t249 VGND 33.717
R720 VGND.t207 VGND.t99 33.717
R721 VGND.n1253 VGND.n1218 33.5064
R722 VGND.n1376 VGND.t196 33.462
R723 VGND.n1376 VGND.t360 33.462
R724 VGND.n21 VGND.t384 33.462
R725 VGND.n21 VGND.t362 33.462
R726 VGND.n42 VGND.t473 33.462
R727 VGND.n42 VGND.t269 33.462
R728 VGND.n1201 VGND.t206 33.462
R729 VGND.n1201 VGND.t406 33.462
R730 VGND.n1199 VGND.t9 33.462
R731 VGND.n1199 VGND.t439 33.462
R732 VGND.n199 VGND.t229 33.462
R733 VGND.n199 VGND.t433 33.462
R734 VGND.n391 VGND.t100 33.462
R735 VGND.n391 VGND.t135 33.462
R736 VGND.n406 VGND.t459 33.462
R737 VGND.n406 VGND.t66 33.462
R738 VGND.n161 VGND.t54 33.462
R739 VGND.n161 VGND.t418 33.462
R740 VGND.n126 VGND.t251 33.462
R741 VGND.n126 VGND.t133 33.462
R742 VGND.n58 VGND.t210 33.462
R743 VGND.n58 VGND.t72 33.462
R744 VGND.n1284 VGND.n1198 30.8711
R745 VGND.n1263 VGND.n1206 30.4946
R746 VGND.n560 VGND.n559 29.66
R747 VGND.n664 VGND.n396 28.9887
R748 VGND.n1251 VGND.t431 28.3801
R749 VGND.n1271 VGND.t461 28.3801
R750 VGND.n1197 VGND.t310 28.3801
R751 VGND.n1231 VGND.t453 28.3166
R752 VGND.n1378 VGND.n1348 28.2358
R753 VGND.n1334 VGND.n16 28.2358
R754 VGND.n281 VGND.n280 28.2358
R755 VGND.n249 VGND.n248 28.2358
R756 VGND.n108 VGND.n74 28.2358
R757 VGND.n220 VGND.n219 26.314
R758 VGND.n1136 VGND.n1135 26.314
R759 VGND.n1278 VGND.n1277 25.977
R760 VGND.n210 VGND.n209 25.977
R761 VGND.n675 VGND.n674 25.977
R762 VGND.n395 VGND.t19 25.9346
R763 VGND.n263 VGND.n256 25.7355
R764 VGND.n268 VGND.n254 25.7355
R765 VGND.n879 VGND.n878 25.7355
R766 VGND.n1289 VGND.n1288 25.6926
R767 VGND.n208 VGND.n205 25.6926
R768 VGND.n1131 VGND.n1130 25.6926
R769 VGND.n1184 VGND.n51 25.6926
R770 VGND.n649 VGND.n648 25.666
R771 VGND.n1044 VGND.n1043 25.666
R772 VGND.n1366 VGND.n1364 25.6005
R773 VGND.n1347 VGND.n2 25.6005
R774 VGND.n1330 VGND.n1329 25.6005
R775 VGND.n1314 VGND.n1313 25.6005
R776 VGND.n276 VGND.n252 25.6005
R777 VGND.n296 VGND.n295 25.6005
R778 VGND.n243 VGND.n242 25.6005
R779 VGND.n1265 VGND.n1263 25.6005
R780 VGND.n107 VGND.n106 25.6005
R781 VGND.n95 VGND.n94 25.6005
R782 VGND VGND.t37 25.2879
R783 VGND.t375 VGND.t306 25.2879
R784 VGND.n1169 VGND.n1168 24.9894
R785 VGND.n629 VGND.t387 24.9236
R786 VGND.n629 VGND.t11 24.9236
R787 VGND.n1024 VGND.t312 24.9236
R788 VGND.n1024 VGND.t437 24.9236
R789 VGND.n1022 VGND.t272 24.9236
R790 VGND.n1022 VGND.t391 24.9236
R791 VGND.n1019 VGND.t398 24.9236
R792 VGND.n1019 VGND.t276 24.9236
R793 VGND.n656 VGND.t314 24.6931
R794 VGND.n1023 VGND.t491 24.6931
R795 VGND.n1010 VGND.t496 24.6931
R796 VGND.n1367 VGND.n1366 24.4711
R797 VGND.n1371 VGND.n1351 24.4711
R798 VGND.n1336 VGND.n2 24.4711
R799 VGND.n1335 VGND.n1334 24.4711
R800 VGND.n1329 VGND.n1328 24.4711
R801 VGND.n1324 VGND.n20 24.4711
R802 VGND.n1313 VGND.n1312 24.4711
R803 VGND.n256 VGND.n29 24.4711
R804 VGND.n273 VGND.n254 24.4711
R805 VGND.n276 VGND.n274 24.4711
R806 VGND.n283 VGND.n281 24.4711
R807 VGND.n295 VGND.n250 24.4711
R808 VGND.n248 VGND.n237 24.4711
R809 VGND.n244 VGND.n243 24.4711
R810 VGND.n106 VGND.n105 24.4711
R811 VGND.n101 VGND.n78 24.4711
R812 VGND.n100 VGND.n80 24.4711
R813 VGND.n96 VGND.n95 24.4711
R814 VGND.n1367 VGND.n1351 24.0946
R815 VGND.n1336 VGND.n1335 24.0946
R816 VGND.n1328 VGND.n20 24.0946
R817 VGND.n1312 VGND.n29 24.0946
R818 VGND.n274 VGND.n273 24.0946
R819 VGND.n283 VGND.n250 24.0946
R820 VGND.n244 VGND.n237 24.0946
R821 VGND.n1253 VGND.n1252 24.0946
R822 VGND.n1273 VGND.n1272 24.0946
R823 VGND.n209 VGND.n208 24.0946
R824 VGND.n105 VGND.n78 24.0946
R825 VGND.n96 VGND.n80 24.0946
R826 VGND.n196 VGND.t499 24.0005
R827 VGND.n203 VGND.t489 24.0005
R828 VGND.n328 VGND.t389 24.0005
R829 VGND.n1319 VGND.n1318 23.7181
R830 VGND.n780 VGND.n183 23.7181
R831 VGND.n780 VGND.n779 23.7181
R832 VGND.n873 VGND.n841 23.7181
R833 VGND.n1189 VGND.n1188 23.7181
R834 VGND.n1247 VGND.n1244 22.9652
R835 VGND.n663 VGND.n662 22.9652
R836 VGND.n1377 VGND.n1349 22.2123
R837 VGND.n1378 VGND.n1377 22.2123
R838 VGND.n1323 VGND.n22 22.2123
R839 VGND.n1319 VGND.n22 22.2123
R840 VGND.n1273 VGND.n1202 22.2123
R841 VGND.n1278 VGND.n1200 22.2123
R842 VGND.n219 VGND.n200 22.2123
R843 VGND.n215 VGND.n200 22.2123
R844 VGND.n878 VGND.n162 22.2123
R845 VGND.n874 VGND.n162 22.2123
R846 VGND.n1135 VGND.n127 22.2123
R847 VGND.n1131 VGND.n127 22.2123
R848 VGND.n1168 VGND.n59 22.2123
R849 VGND.n74 VGND.n59 22.2123
R850 VGND.n627 VGND.t428 22.0959
R851 VGND.n393 VGND.t208 22.0959
R852 VGND.n568 VGND.t475 21.795
R853 VGND.n1247 VGND.n1219 21.4593
R854 VGND.n1284 VGND.n1283 21.4593
R855 VGND.n662 VGND.n626 21.4593
R856 VGND.n674 VGND.n396 21.4593
R857 VGND.n1052 VGND.n1051 21.0829
R858 VGND.n1058 VGND.n1057 20.6669
R859 VGND.n1364 VGND.n1353 19.9534
R860 VGND.n1348 VGND.n1347 19.9534
R861 VGND.n1330 VGND.n16 19.9534
R862 VGND.n1314 VGND.n23 19.9534
R863 VGND.n280 VGND.n252 19.9534
R864 VGND.n296 VGND.n249 19.9534
R865 VGND.n242 VGND.n163 19.9534
R866 VGND.n1244 VGND.n1243 19.9534
R867 VGND.n108 VGND.n107 19.9534
R868 VGND.n94 VGND.n83 19.9534
R869 VGND.n1243 VGND.n1222 19.577
R870 VGND.n1360 VGND.n1353 19.3355
R871 VGND.n90 VGND.n83 19.3355
R872 VGND.n561 VGND.n558 19.0176
R873 VGND.n651 VGND.n630 18.824
R874 VGND.n1046 VGND.n1025 18.824
R875 VGND.n335 VGND.n330 18.2791
R876 VGND.n1082 VGND.n1081 18.2791
R877 VGND.n1318 VGND.n23 17.3181
R878 VGND.n834 VGND.n163 17.3181
R879 VGND.n1230 VGND.n1229 17.3181
R880 VGND.n541 VGND.n540 17.2917
R881 VGND.n592 VGND.n591 17.1022
R882 VGND.n849 VGND.n848 16.9545
R883 VGND.n1252 VGND.n1219 16.9417
R884 VGND.t268 VGND.t303 16.8587
R885 VGND.t440 VGND.t430 16.8587
R886 VGND.t234 VGND.t43 16.8587
R887 VGND.t434 VGND.t230 16.8587
R888 VGND.t153 VGND.t474 16.8587
R889 VGND.t123 VGND.t415 16.8587
R890 VGND.n826 VGND.n167 16.7924
R891 VGND.n917 VGND.n916 16.4139
R892 VGND.n561 VGND.n560 16.217
R893 VGND.n654 VGND.n630 15.8123
R894 VGND.n1049 VGND.n1025 15.8123
R895 VGND.n552 VGND.n412 15.5279
R896 VGND.n1057 VGND.n1020 15.4358
R897 VGND.n640 VGND.n639 14.8179
R898 VGND.n1035 VGND.n1034 14.8179
R899 VGND.n784 VGND.n183 14.775
R900 VGND.n796 VGND.n792 14.775
R901 VGND.n360 VGND.n359 14.775
R902 VGND.n869 VGND.n841 14.775
R903 VGND.n1189 VGND.n49 14.775
R904 VGND.n834 VGND.n833 14.775
R905 VGND.n680 VGND.n679 14.6434
R906 VGND.n436 VGND.n418 13.8859
R907 VGND.n907 VGND.n148 13.8859
R908 VGND.n1239 VGND.n1222 13.5534
R909 VGND.n549 VGND.n412 13.177
R910 VGND.n1267 VGND.n1265 12.8005
R911 VGND.n583 VGND.n578 12.8005
R912 VGND.n1051 VGND.n1050 12.8005
R913 VGND.n512 VGND.n466 12.3514
R914 VGND.n540 VGND.n448 12.3514
R915 VGND.n513 VGND.n512 12.1268
R916 VGND.n1237 VGND.n1224 12.0476
R917 VGND.n1239 VGND.n1237 11.6711
R918 VGND.n1277 VGND.n1202 11.2946
R919 VGND.n675 VGND.n392 11.2946
R920 VGND.n1267 VGND.n1204 10.9181
R921 VGND.n779 VGND.n184 10.5983
R922 VGND.n1283 VGND.n1200 10.5417
R923 VGND.n1232 VGND.n1230 9.78874
R924 VGND.n1356 VGND.n1355 9.71789
R925 VGND.n159 VGND.n158 9.71789
R926 VGND.n86 VGND.n85 9.71789
R927 VGND.n819 VGND.n818 9.71789
R928 VGND.n658 VGND.n657 9.41227
R929 VGND.n206 VGND.n205 9.3005
R930 VGND.n1298 VGND.n1297 9.3005
R931 VGND.n1296 VGND.n1295 9.3005
R932 VGND.n1290 VGND.n1289 9.3005
R933 VGND.n1286 VGND.n1196 9.3005
R934 VGND.n1283 VGND.n1281 9.3005
R935 VGND.n1277 VGND.n1276 9.3005
R936 VGND.n1272 VGND.n1270 9.3005
R937 VGND.n1268 VGND.n1267 9.3005
R938 VGND.n1217 VGND.n1208 9.3005
R939 VGND.n1252 VGND.n1250 9.3005
R940 VGND.n1248 VGND.n1247 9.3005
R941 VGND.n1241 VGND.n1222 9.3005
R942 VGND.n1237 VGND.n1235 9.3005
R943 VGND.n1233 VGND.n1232 9.3005
R944 VGND.n1230 VGND.n1225 9.3005
R945 VGND.n1234 VGND.n1224 9.3005
R946 VGND.n1240 VGND.n1239 9.3005
R947 VGND.n1243 VGND.n1242 9.3005
R948 VGND.n1244 VGND.n1221 9.3005
R949 VGND.n1249 VGND.n1219 9.3005
R950 VGND.n1254 VGND.n1253 9.3005
R951 VGND.n1263 VGND.n1262 9.3005
R952 VGND.n1265 VGND.n1205 9.3005
R953 VGND.n1269 VGND.n1204 9.3005
R954 VGND.n1274 VGND.n1273 9.3005
R955 VGND.n1275 VGND.n1202 9.3005
R956 VGND.n1279 VGND.n1278 9.3005
R957 VGND.n1280 VGND.n1200 9.3005
R958 VGND.n1285 VGND.n1284 9.3005
R959 VGND.n1288 VGND.n1287 9.3005
R960 VGND.n208 VGND.n207 9.3005
R961 VGND.n209 VGND.n202 9.3005
R962 VGND.n211 VGND.n210 9.3005
R963 VGND.n212 VGND.n201 9.3005
R964 VGND.n214 VGND.n213 9.3005
R965 VGND.n216 VGND.n215 9.3005
R966 VGND.n217 VGND.n200 9.3005
R967 VGND.n219 VGND.n218 9.3005
R968 VGND.n221 VGND.n220 9.3005
R969 VGND.n223 VGND.n222 9.3005
R970 VGND.n224 VGND.n194 9.3005
R971 VGND.n226 VGND.n225 9.3005
R972 VGND.n227 VGND.n191 9.3005
R973 VGND.n764 VGND.n763 9.3005
R974 VGND.n753 VGND.n189 9.3005
R975 VGND.n770 VGND.n769 9.3005
R976 VGND.n771 VGND.n186 9.3005
R977 VGND.n773 VGND.n772 9.3005
R978 VGND.n774 VGND.n185 9.3005
R979 VGND.n777 VGND.n776 9.3005
R980 VGND.n796 VGND.n795 9.3005
R981 VGND.n792 VGND.n791 9.3005
R982 VGND.n790 VGND.n789 9.3005
R983 VGND.n788 VGND.n178 9.3005
R984 VGND.n784 VGND.n783 9.3005
R985 VGND.n782 VGND.n183 9.3005
R986 VGND.n781 VGND.n780 9.3005
R987 VGND.n779 VGND.n778 9.3005
R988 VGND.n713 VGND.n712 9.3005
R989 VGND.n715 VGND.n714 9.3005
R990 VGND.n716 VGND.n316 9.3005
R991 VGND.n718 VGND.n717 9.3005
R992 VGND.n719 VGND.n315 9.3005
R993 VGND.n721 VGND.n720 9.3005
R994 VGND.n722 VGND.n314 9.3005
R995 VGND.n724 VGND.n723 9.3005
R996 VGND.n726 VGND.n725 9.3005
R997 VGND.n711 VGND.n710 9.3005
R998 VGND.n709 VGND.n320 9.3005
R999 VGND.n331 VGND.n330 9.3005
R1000 VGND.n335 VGND.n334 9.3005
R1001 VGND.n700 VGND.n699 9.3005
R1002 VGND.n698 VGND.n327 9.3005
R1003 VGND.n697 VGND.n696 9.3005
R1004 VGND.n695 VGND.n385 9.3005
R1005 VGND.n694 VGND.n693 9.3005
R1006 VGND.n690 VGND.n386 9.3005
R1007 VGND.n688 VGND.n687 9.3005
R1008 VGND.n686 VGND.n685 9.3005
R1009 VGND.n684 VGND.n389 9.3005
R1010 VGND.n683 VGND.n682 9.3005
R1011 VGND.n681 VGND.n680 9.3005
R1012 VGND.n677 VGND.n392 9.3005
R1013 VGND.n647 VGND.n646 9.3005
R1014 VGND.n645 VGND.n644 9.3005
R1015 VGND.n640 VGND.n635 9.3005
R1016 VGND.n649 VGND.n631 9.3005
R1017 VGND.n652 VGND.n651 9.3005
R1018 VGND.n654 VGND.n653 9.3005
R1019 VGND.n655 VGND.n628 9.3005
R1020 VGND.n659 VGND.n658 9.3005
R1021 VGND.n660 VGND.n626 9.3005
R1022 VGND.n662 VGND.n661 9.3005
R1023 VGND.n663 VGND.n625 9.3005
R1024 VGND.n665 VGND.n664 9.3005
R1025 VGND.n398 VGND.n396 9.3005
R1026 VGND.n674 VGND.n673 9.3005
R1027 VGND.n676 VGND.n675 9.3005
R1028 VGND.n679 VGND.n678 9.3005
R1029 VGND.n727 VGND.n311 9.3005
R1030 VGND.n730 VGND.n729 9.3005
R1031 VGND.n731 VGND.n310 9.3005
R1032 VGND.n359 VGND.n357 9.3005
R1033 VGND.n360 VGND.n341 9.3005
R1034 VGND.n365 VGND.n364 9.3005
R1035 VGND.n382 VGND.n381 9.3005
R1036 VGND.n380 VGND.n339 9.3005
R1037 VGND.n379 VGND.n378 9.3005
R1038 VGND.n377 VGND.n367 9.3005
R1039 VGND.n376 VGND.n375 9.3005
R1040 VGND.n374 VGND.n369 9.3005
R1041 VGND.n373 VGND.n372 9.3005
R1042 VGND.n370 VGND.n309 9.3005
R1043 VGND.n744 VGND.n743 9.3005
R1044 VGND.n740 VGND.n739 9.3005
R1045 VGND.n591 VGND.n590 9.3005
R1046 VGND.n589 VGND.n588 9.3005
R1047 VGND.n586 VGND.n574 9.3005
R1048 VGND.n593 VGND.n572 9.3005
R1049 VGND.n596 VGND.n595 9.3005
R1050 VGND.n597 VGND.n571 9.3005
R1051 VGND.n599 VGND.n598 9.3005
R1052 VGND.n601 VGND.n570 9.3005
R1053 VGND.n603 VGND.n602 9.3005
R1054 VGND.n612 VGND.n611 9.3005
R1055 VGND.n614 VGND.n613 9.3005
R1056 VGND.n567 VGND.n566 9.3005
R1057 VGND.n565 VGND.n407 9.3005
R1058 VGND.n426 VGND.n418 9.3005
R1059 VGND.n436 VGND.n435 9.3005
R1060 VGND.n438 VGND.n415 9.3005
R1061 VGND.n442 VGND.n441 9.3005
R1062 VGND.n443 VGND.n414 9.3005
R1063 VGND.n546 VGND.n444 9.3005
R1064 VGND.n545 VGND.n544 9.3005
R1065 VGND.n543 VGND.n542 9.3005
R1066 VGND.n540 VGND.n539 9.3005
R1067 VGND.n538 VGND.n537 9.3005
R1068 VGND.n535 VGND.n449 9.3005
R1069 VGND.n534 VGND.n533 9.3005
R1070 VGND.n532 VGND.n450 9.3005
R1071 VGND.n459 VGND.n458 9.3005
R1072 VGND.n463 VGND.n462 9.3005
R1073 VGND.n523 VGND.n522 9.3005
R1074 VGND.n520 VGND.n457 9.3005
R1075 VGND.n518 VGND.n517 9.3005
R1076 VGND.n516 VGND.n464 9.3005
R1077 VGND.n515 VGND.n514 9.3005
R1078 VGND.n512 VGND.n511 9.3005
R1079 VGND.n510 VGND.n509 9.3005
R1080 VGND.n507 VGND.n467 9.3005
R1081 VGND.n506 VGND.n505 9.3005
R1082 VGND.n504 VGND.n468 9.3005
R1083 VGND.n503 VGND.n502 9.3005
R1084 VGND.n501 VGND.n469 9.3005
R1085 VGND.n500 VGND.n499 9.3005
R1086 VGND.n498 VGND.n497 9.3005
R1087 VGND.n495 VGND.n494 9.3005
R1088 VGND.n474 VGND.n472 9.3005
R1089 VGND.n486 VGND.n485 9.3005
R1090 VGND.n482 VGND.n413 9.3005
R1091 VGND.n550 VGND.n549 9.3005
R1092 VGND.n551 VGND.n412 9.3005
R1093 VGND.n552 VGND 9.3005
R1094 VGND.n555 VGND.n554 9.3005
R1095 VGND.n88 VGND.n84 9.3005
R1096 VGND.n91 VGND.n90 9.3005
R1097 VGND.n92 VGND.n83 9.3005
R1098 VGND.n94 VGND.n93 9.3005
R1099 VGND.n95 VGND.n81 9.3005
R1100 VGND.n97 VGND.n96 9.3005
R1101 VGND.n98 VGND.n80 9.3005
R1102 VGND.n100 VGND.n99 9.3005
R1103 VGND.n102 VGND.n101 9.3005
R1104 VGND.n103 VGND.n78 9.3005
R1105 VGND.n105 VGND.n104 9.3005
R1106 VGND.n106 VGND.n76 9.3005
R1107 VGND.n107 VGND.n66 9.3005
R1108 VGND.n109 VGND.n108 9.3005
R1109 VGND.n74 VGND.n73 9.3005
R1110 VGND.n67 VGND.n59 9.3005
R1111 VGND.n1168 VGND.n1167 9.3005
R1112 VGND.n1170 VGND.n1169 9.3005
R1113 VGND.n1172 VGND.n1171 9.3005
R1114 VGND.n55 VGND.n54 9.3005
R1115 VGND.n1178 VGND.n1177 9.3005
R1116 VGND.n1179 VGND.n53 9.3005
R1117 VGND.n1181 VGND.n1180 9.3005
R1118 VGND.n1182 VGND.n52 9.3005
R1119 VGND.n1185 VGND.n1184 9.3005
R1120 VGND.n1186 VGND.n51 9.3005
R1121 VGND.n1188 VGND.n1187 9.3005
R1122 VGND.n1189 VGND.n50 9.3005
R1123 VGND.n1116 VGND.n49 9.3005
R1124 VGND.n1121 VGND.n1120 9.3005
R1125 VGND.n1117 VGND.n131 9.3005
R1126 VGND.n1130 VGND.n1129 9.3005
R1127 VGND.n1132 VGND.n1131 9.3005
R1128 VGND.n1133 VGND.n127 9.3005
R1129 VGND.n1135 VGND.n1134 9.3005
R1130 VGND.n1137 VGND.n1136 9.3005
R1131 VGND.n1139 VGND.n1138 9.3005
R1132 VGND.n1140 VGND.n124 9.3005
R1133 VGND.n1142 VGND.n1141 9.3005
R1134 VGND.n1144 VGND.n1143 9.3005
R1135 VGND.n1145 VGND.n122 9.3005
R1136 VGND.n1147 VGND.n1146 9.3005
R1137 VGND.n1148 VGND.n121 9.3005
R1138 VGND.n1150 VGND.n1149 9.3005
R1139 VGND.n1151 VGND.n119 9.3005
R1140 VGND.n1153 VGND.n1152 9.3005
R1141 VGND.n848 VGND.n118 9.3005
R1142 VGND.n882 VGND.n881 9.3005
R1143 VGND.n879 VGND.n157 9.3005
R1144 VGND.n878 VGND.n877 9.3005
R1145 VGND.n876 VGND.n162 9.3005
R1146 VGND.n875 VGND.n874 9.3005
R1147 VGND.n873 VGND.n872 9.3005
R1148 VGND.n871 VGND.n841 9.3005
R1149 VGND.n870 VGND.n869 9.3005
R1150 VGND.n867 VGND.n842 9.3005
R1151 VGND.n866 VGND.n865 9.3005
R1152 VGND.n864 VGND.n843 9.3005
R1153 VGND.n863 VGND.n862 9.3005
R1154 VGND.n845 VGND.n844 9.3005
R1155 VGND.n857 VGND.n856 9.3005
R1156 VGND.n850 VGND.n849 9.3005
R1157 VGND.n1054 VGND.n1053 9.3005
R1158 VGND.n1047 VGND.n1046 9.3005
R1159 VGND.n1042 VGND.n1041 9.3005
R1160 VGND.n1035 VGND.n1030 9.3005
R1161 VGND.n1040 VGND.n1039 9.3005
R1162 VGND.n1044 VGND.n1026 9.3005
R1163 VGND.n1049 VGND.n1048 9.3005
R1164 VGND.n1050 VGND.n1021 9.3005
R1165 VGND.n1055 VGND.n1020 9.3005
R1166 VGND.n894 VGND.n148 9.3005
R1167 VGND.n907 VGND.n906 9.3005
R1168 VGND.n909 VGND.n145 9.3005
R1169 VGND.n913 VGND.n912 9.3005
R1170 VGND.n914 VGND.n144 9.3005
R1171 VGND.n1057 VGND.n1056 9.3005
R1172 VGND.n1081 VGND.n1080 9.3005
R1173 VGND VGND.n1079 9.3005
R1174 VGND.n1078 VGND.n1077 9.3005
R1175 VGND.n1076 VGND.n998 9.3005
R1176 VGND.n1075 VGND.n1074 9.3005
R1177 VGND.n1073 VGND.n999 9.3005
R1178 VGND.n1072 VGND 9.3005
R1179 VGND.n1071 VGND.n1002 9.3005
R1180 VGND.n1014 VGND.n1013 9.3005
R1181 VGND.n1018 VGND.n1017 9.3005
R1182 VGND.n1062 VGND.n1061 9.3005
R1183 VGND.n1058 VGND.n1009 9.3005
R1184 VGND.n1089 VGND.n1088 9.3005
R1185 VGND.n1087 VGND.n994 9.3005
R1186 VGND.n1086 VGND.n1085 9.3005
R1187 VGND.n1082 VGND.n995 9.3005
R1188 VGND.n1092 VGND.n1091 9.3005
R1189 VGND.n1093 VGND.n142 9.3005
R1190 VGND.n1102 VGND.n1101 9.3005
R1191 VGND.n1104 VGND.n1103 9.3005
R1192 VGND.n944 VGND.n943 9.3005
R1193 VGND.n945 VGND.n941 9.3005
R1194 VGND.n947 VGND.n946 9.3005
R1195 VGND.n948 VGND.n940 9.3005
R1196 VGND.n950 VGND.n949 9.3005
R1197 VGND.n952 VGND.n939 9.3005
R1198 VGND.n954 VGND.n953 9.3005
R1199 VGND.n956 VGND.n955 9.3005
R1200 VGND.n926 VGND.n921 9.3005
R1201 VGND.n969 VGND.n968 9.3005
R1202 VGND.n967 VGND.n966 9.3005
R1203 VGND.n965 VGND.n929 9.3005
R1204 VGND.n964 VGND.n963 9.3005
R1205 VGND.n962 VGND.n935 9.3005
R1206 VGND.n961 VGND.n960 9.3005
R1207 VGND.n959 VGND.n958 9.3005
R1208 VGND.n984 VGND.n983 9.3005
R1209 VGND.n982 VGND.n981 9.3005
R1210 VGND.n980 VGND.n920 9.3005
R1211 VGND.n978 VGND.n977 9.3005
R1212 VGND.n991 VGND.n915 9.3005
R1213 VGND.n989 VGND.n988 9.3005
R1214 VGND.n823 VGND.n822 9.3005
R1215 VGND.n824 VGND.n167 9.3005
R1216 VGND.n826 VGND.n825 9.3005
R1217 VGND.n828 VGND.n166 9.3005
R1218 VGND.n831 VGND.n830 9.3005
R1219 VGND.n833 VGND.n832 9.3005
R1220 VGND.n834 VGND.n164 9.3005
R1221 VGND.n240 VGND.n163 9.3005
R1222 VGND.n242 VGND.n241 9.3005
R1223 VGND.n243 VGND.n238 9.3005
R1224 VGND.n245 VGND.n244 9.3005
R1225 VGND.n246 VGND.n237 9.3005
R1226 VGND.n248 VGND.n247 9.3005
R1227 VGND.n249 VGND.n235 9.3005
R1228 VGND.n297 VGND.n296 9.3005
R1229 VGND.n295 VGND.n293 9.3005
R1230 VGND.n285 VGND.n250 9.3005
R1231 VGND.n284 VGND.n283 9.3005
R1232 VGND.n281 VGND.n251 9.3005
R1233 VGND.n280 VGND.n279 9.3005
R1234 VGND.n278 VGND.n252 9.3005
R1235 VGND.n277 VGND.n276 9.3005
R1236 VGND.n274 VGND.n253 9.3005
R1237 VGND.n273 VGND.n271 9.3005
R1238 VGND.n270 VGND.n254 9.3005
R1239 VGND.n269 VGND.n268 9.3005
R1240 VGND.n266 VGND.n255 9.3005
R1241 VGND.n263 VGND.n262 9.3005
R1242 VGND.n261 VGND.n256 9.3005
R1243 VGND.n260 VGND.n29 9.3005
R1244 VGND.n1312 VGND.n1311 9.3005
R1245 VGND.n1313 VGND.n26 9.3005
R1246 VGND.n1315 VGND.n1314 9.3005
R1247 VGND.n1316 VGND.n23 9.3005
R1248 VGND.n1318 VGND.n1317 9.3005
R1249 VGND.n1320 VGND.n1319 9.3005
R1250 VGND.n1321 VGND.n22 9.3005
R1251 VGND.n1323 VGND.n1322 9.3005
R1252 VGND.n1325 VGND.n1324 9.3005
R1253 VGND.n1326 VGND.n20 9.3005
R1254 VGND.n1328 VGND.n1327 9.3005
R1255 VGND.n1329 VGND.n17 9.3005
R1256 VGND.n1331 VGND.n1330 9.3005
R1257 VGND.n1332 VGND.n16 9.3005
R1258 VGND.n1334 VGND.n1333 9.3005
R1259 VGND.n1335 VGND.n14 9.3005
R1260 VGND.n1337 VGND.n1336 9.3005
R1261 VGND.n10 VGND.n2 9.3005
R1262 VGND.n1347 VGND.n1346 9.3005
R1263 VGND.n1348 VGND.n0 9.3005
R1264 VGND.n1379 VGND.n1378 9.3005
R1265 VGND.n1377 VGND.n1375 9.3005
R1266 VGND.n1374 VGND.n1349 9.3005
R1267 VGND.n1373 VGND.n1372 9.3005
R1268 VGND.n1371 VGND.n1370 9.3005
R1269 VGND.n1369 VGND.n1351 9.3005
R1270 VGND.n1368 VGND.n1367 9.3005
R1271 VGND.n1366 VGND.n1352 9.3005
R1272 VGND.n1364 VGND.n1363 9.3005
R1273 VGND.n1362 VGND.n1353 9.3005
R1274 VGND.n1361 VGND.n1360 9.3005
R1275 VGND.n1358 VGND.n1354 9.3005
R1276 VGND.n679 VGND.n392 9.03579
R1277 VGND.n549 VGND.n413 9.03579
R1278 VGND VGND.t403 8.42962
R1279 VGND.n204 VGND.n201 8.28285
R1280 VGND.n225 VGND.n224 8.23546
R1281 VGND.n224 VGND.n223 8.23546
R1282 VGND.n685 VGND.n684 8.23546
R1283 VGND.n684 VGND.n683 8.23546
R1284 VGND.n699 VGND.n698 8.23546
R1285 VGND.n698 VGND.n697 8.23546
R1286 VGND.n711 VGND.n320 8.23546
R1287 VGND.n567 VGND.n407 8.23546
R1288 VGND.n613 VGND.n567 8.23546
R1289 VGND.n613 VGND.n612 8.23546
R1290 VGND.n602 VGND.n601 8.23546
R1291 VGND.n599 VGND.n571 8.23546
R1292 VGND.n595 VGND.n571 8.23546
R1293 VGND.n1152 VGND.n1151 8.23546
R1294 VGND.n1151 VGND.n1150 8.23546
R1295 VGND.n1150 VGND.n121 8.23546
R1296 VGND.n1146 VGND.n121 8.23546
R1297 VGND.n1146 VGND.n1145 8.23546
R1298 VGND.n1145 VGND.n1144 8.23546
R1299 VGND.n1141 VGND.n1140 8.23546
R1300 VGND.n1140 VGND.n1139 8.23546
R1301 VGND.n1079 VGND.n1078 8.23546
R1302 VGND.n1078 VGND.n998 8.23546
R1303 VGND.n1074 VGND.n1073 8.23546
R1304 VGND.n1073 VGND.n1072 8.23546
R1305 VGND.n1072 VGND.n1002 8.23546
R1306 VGND.n1061 VGND.n1018 8.23546
R1307 VGND.n1089 VGND.n994 8.23546
R1308 VGND.n1085 VGND.n994 8.23546
R1309 VGND.n563 VGND.n562 8.16157
R1310 VGND.n612 VGND.n569 8.05644
R1311 VGND.n683 VGND.n390 7.6984
R1312 VGND.n329 VGND.n320 7.6984
R1313 VGND.n595 VGND.n594 7.6984
R1314 VGND.n1152 VGND.n120 7.6984
R1315 VGND.n1139 VGND.n125 7.6984
R1316 VGND.n1079 VGND.n997 7.6984
R1317 VGND.n1074 VGND.n1000 7.6984
R1318 VGND.n484 VGND.n413 7.51354
R1319 VGND.n1084 VGND.n1083 7.16134
R1320 VGND.n1232 VGND.n1224 7.15344
R1321 VGND.n382 VGND.n339 7.15139
R1322 VGND.n712 VGND.n711 7.11268
R1323 VGND.n697 VGND.n385 6.90655
R1324 VGND.n1272 VGND.n1204 6.77697
R1325 VGND.n690 VGND.n689 6.63802
R1326 VGND.n363 VGND.n340 6.61527
R1327 VGND.n986 VGND.n918 6.57117
R1328 VGND.n986 VGND.n985 6.57117
R1329 VGND.n764 VGND.n191 6.56535
R1330 VGND.n789 VGND.n788 6.26433
R1331 VGND.n1297 VGND.n1296 6.26433
R1332 VGND.n546 VGND.n545 6.26433
R1333 VGND.n867 VGND.n866 6.26433
R1334 VGND.n866 VGND.n843 6.26433
R1335 VGND.n1120 VGND.n1117 6.26433
R1336 VGND.n1182 VGND.n1181 6.26433
R1337 VGND.n1181 VGND.n53 6.26433
R1338 VGND.n830 VGND.n828 6.26433
R1339 VGND.n587 VGND.n586 6.19624
R1340 VGND.n740 VGND.n310 6.02861
R1341 VGND.n727 VGND.n726 6.02861
R1342 VGND.n950 VGND.n940 6.0286
R1343 VGND.n1359 VGND.n1358 5.98311
R1344 VGND.n267 VGND.n266 5.98311
R1345 VGND.n644 VGND.n634 5.98311
R1346 VGND.n881 VGND.n880 5.98311
R1347 VGND.n89 VGND.n88 5.98311
R1348 VGND.n1039 VGND.n1029 5.98311
R1349 VGND.n822 VGND.n821 5.98311
R1350 VGND.n1297 VGND.n43 5.85582
R1351 VGND.n364 VGND.n361 5.85582
R1352 VGND.n554 VGND.n553 5.85582
R1353 VGND.n588 VGND.n573 5.85582
R1354 VGND.n868 VGND.n867 5.85582
R1355 VGND.n1117 VGND.n129 5.85582
R1356 VGND.n1183 VGND.n1182 5.85582
R1357 VGND.n828 VGND.n827 5.85582
R1358 VGND.n978 VGND.n921 5.80542
R1359 VGND.n862 VGND.n843 5.65809
R1360 VGND.n1177 VGND.n53 5.65809
R1361 VGND.n382 VGND.n338 5.63966
R1362 VGND.n408 VGND.n407 5.63966
R1363 VGND.n789 VGND.n179 5.51539
R1364 VGND.n546 VGND.n414 5.37524
R1365 VGND.n991 VGND.n144 5.37524
R1366 VGND.n990 VGND.n916 5.29405
R1367 VGND.n1013 VGND.n1011 5.19211
R1368 VGND.n796 VGND.n793 5.13108
R1369 VGND.n796 VGND.n794 5.13108
R1370 VGND.n1229 VGND.n1226 5.13108
R1371 VGND.n1229 VGND.n1228 5.13108
R1372 VGND.n639 VGND.n636 5.13108
R1373 VGND.n639 VGND.n638 5.13108
R1374 VGND.n359 VGND.n342 5.13108
R1375 VGND.n359 VGND.n358 5.13108
R1376 VGND.n578 VGND.n576 5.13108
R1377 VGND.n578 VGND.n577 5.13108
R1378 VGND.n418 VGND.n416 5.13108
R1379 VGND.n418 VGND.n417 5.13108
R1380 VGND.n148 VGND.n146 5.13108
R1381 VGND.n148 VGND.n147 5.13108
R1382 VGND.n1034 VGND.n1031 5.13108
R1383 VGND.n1034 VGND.n1033 5.13108
R1384 VGND.n223 VGND.n197 4.92358
R1385 VGND.n542 VGND.n445 4.90263
R1386 VGND.n767 VGND.n190 4.85762
R1387 VGND.n1175 VGND.n1174 4.85762
R1388 VGND.n860 VGND.n859 4.85762
R1389 VGND.n1358 VGND.n1357 4.8005
R1390 VGND.n266 VGND.n265 4.8005
R1391 VGND.n644 VGND.n643 4.8005
R1392 VGND.n881 VGND.n160 4.8005
R1393 VGND.n88 VGND.n87 4.8005
R1394 VGND.n1039 VGND.n1038 4.8005
R1395 VGND.n822 VGND.n820 4.8005
R1396 VGND.n378 VGND.n377 4.67352
R1397 VGND.n377 VGND.n376 4.67352
R1398 VGND.n376 VGND.n369 4.67352
R1399 VGND.n372 VGND.n309 4.67352
R1400 VGND.n743 VGND.n309 4.67352
R1401 VGND.n723 VGND.n722 4.67352
R1402 VGND.n722 VGND.n721 4.67352
R1403 VGND.n721 VGND.n315 4.67352
R1404 VGND.n717 VGND.n716 4.67352
R1405 VGND.n716 VGND.n715 4.67352
R1406 VGND.n507 VGND.n506 4.67352
R1407 VGND.n506 VGND.n468 4.67352
R1408 VGND.n502 VGND.n468 4.67352
R1409 VGND.n502 VGND.n501 4.67352
R1410 VGND.n501 VGND.n500 4.67352
R1411 VGND.n495 VGND.n472 4.67352
R1412 VGND.n535 VGND.n534 4.67352
R1413 VGND.n534 VGND.n450 4.67352
R1414 VGND.n458 VGND.n450 4.67352
R1415 VGND.n463 VGND.n458 4.67352
R1416 VGND.n522 VGND.n463 4.67352
R1417 VGND.n518 VGND.n464 4.67352
R1418 VGND.n946 VGND.n945 4.67352
R1419 VGND.n945 VGND.n944 4.67352
R1420 VGND.n1103 VGND.n1102 4.67352
R1421 VGND.n1102 VGND.n142 4.67352
R1422 VGND.n953 VGND.n952 4.67352
R1423 VGND.n968 VGND.n967 4.67352
R1424 VGND.n967 VGND.n929 4.67352
R1425 VGND.n963 VGND.n962 4.67352
R1426 VGND.n962 VGND.n961 4.67352
R1427 VGND.n340 VGND.n338 4.63943
R1428 VGND.n563 VGND.n408 4.63943
R1429 VGND.n797 VGND.n796 4.62124
R1430 VGND.n359 VGND.n343 4.62124
R1431 VGND.n434 VGND.n418 4.62124
R1432 VGND.n905 VGND.n148 4.62124
R1433 VGND.n366 VGND.n340 4.62124
R1434 VGND.n564 VGND.n563 4.62124
R1435 VGND.n987 VGND.n986 4.62124
R1436 VGND.n514 VGND.n513 4.60638
R1437 VGND.n509 VGND.n466 4.55559
R1438 VGND.n537 VGND.n448 4.55559
R1439 VGND.n300 VGND.n232 4.51401
R1440 VGND.n290 VGND.n286 4.51401
R1441 VGND.n1340 VGND.n8 4.51401
R1442 VGND.n1345 VGND.n1344 4.51401
R1443 VGND.n1070 VGND.n1069 4.51401
R1444 VGND.n1064 VGND.n1063 4.51401
R1445 VGND.n531 VGND.n530 4.51401
R1446 VGND.n525 VGND.n524 4.51401
R1447 VGND.n815 VGND.n168 4.51401
R1448 VGND.n1213 VGND.n1211 4.51401
R1449 VGND.n1256 VGND.n1255 4.51401
R1450 VGND.n1301 VGND.n39 4.51401
R1451 VGND.n1292 VGND.n1291 4.51401
R1452 VGND.n756 VGND.n187 4.51401
R1453 VGND.n760 VGND.n228 4.51401
R1454 VGND.n798 VGND.n176 4.51401
R1455 VGND.n621 VGND.n394 4.51401
R1456 VGND.n667 VGND.n666 4.51401
R1457 VGND.n708 VGND.n707 4.51401
R1458 VGND.n702 VGND.n701 4.51401
R1459 VGND.n747 VGND.n306 4.51401
R1460 VGND.n736 VGND.n732 4.51401
R1461 VGND.n354 VGND.n345 4.51401
R1462 VGND.n904 VGND.n903 4.51401
R1463 VGND.n883 VGND.n156 4.51401
R1464 VGND.n433 VGND.n432 4.51401
R1465 VGND.n617 VGND.n404 4.51401
R1466 VGND.n608 VGND.n604 4.51401
R1467 VGND.n478 VGND.n471 4.51401
R1468 VGND.n488 VGND.n487 4.51401
R1469 VGND.n1107 VGND.n138 4.51401
R1470 VGND.n1098 VGND.n1094 4.51401
R1471 VGND.n1112 VGND.n128 4.51401
R1472 VGND.n1123 VGND.n1122 4.51401
R1473 VGND.n855 VGND.n854 4.51401
R1474 VGND.n1154 VGND.n115 4.51401
R1475 VGND.n1166 VGND.n1165 4.51401
R1476 VGND.n111 VGND.n110 4.51401
R1477 VGND.n976 VGND.n975 4.51401
R1478 VGND.n934 VGND.n933 4.51401
R1479 VGND.n259 VGND.n258 4.51401
R1480 VGND.n1305 VGND.n25 4.51401
R1481 VGND.n755 VGND.n754 4.5005
R1482 VGND.n751 VGND.n192 4.5005
R1483 VGND.n762 VGND.n761 4.5005
R1484 VGND.n1300 VGND.n1299 4.5005
R1485 VGND.n45 VGND.n41 4.5005
R1486 VGND.n1294 VGND.n1293 4.5005
R1487 VGND.n1212 VGND.n1207 4.5005
R1488 VGND.n1261 VGND.n1260 4.5005
R1489 VGND.n1216 VGND.n1210 4.5005
R1490 VGND.n803 VGND.n175 4.5005
R1491 VGND.n800 VGND.n799 4.5005
R1492 VGND.n322 VGND.n321 4.5005
R1493 VGND.n333 VGND.n332 4.5005
R1494 VGND.n326 VGND.n325 4.5005
R1495 VGND.n620 VGND.n397 4.5005
R1496 VGND.n672 VGND.n671 4.5005
R1497 VGND.n624 VGND.n400 4.5005
R1498 VGND.n746 VGND.n745 4.5005
R1499 VGND.n733 VGND.n308 4.5005
R1500 VGND.n738 VGND.n737 4.5005
R1501 VGND.n347 VGND.n344 4.5005
R1502 VGND.n356 VGND.n355 4.5005
R1503 VGND.n616 VGND.n615 4.5005
R1504 VGND.n605 VGND 4.5005
R1505 VGND.n610 VGND.n609 4.5005
R1506 VGND.n428 VGND.n427 4.5005
R1507 VGND.n420 VGND.n419 4.5005
R1508 VGND.n452 VGND.n451 4.5005
R1509 VGND.n461 VGND.n460 4.5005
R1510 VGND.n456 VGND.n455 4.5005
R1511 VGND.n477 VGND.n473 4.5005
R1512 VGND.n493 VGND.n492 4.5005
R1513 VGND.n481 VGND.n476 4.5005
R1514 VGND.n853 VGND.n851 4.5005
R1515 VGND VGND.n117 4.5005
R1516 VGND.n1156 VGND.n1155 4.5005
R1517 VGND.n1111 VGND.n130 4.5005
R1518 VGND.n1128 VGND.n1127 4.5005
R1519 VGND.n1115 VGND.n133 4.5005
R1520 VGND.n888 VGND.n155 4.5005
R1521 VGND.n885 VGND.n884 4.5005
R1522 VGND.n61 VGND.n60 4.5005
R1523 VGND.n71 VGND.n70 4.5005
R1524 VGND.n72 VGND.n65 4.5005
R1525 VGND.n1106 VGND.n1105 4.5005
R1526 VGND.n1095 VGND.n140 4.5005
R1527 VGND.n1100 VGND.n1099 4.5005
R1528 VGND.n1004 VGND.n1003 4.5005
R1529 VGND.n1016 VGND.n1015 4.5005
R1530 VGND.n1008 VGND.n1007 4.5005
R1531 VGND.n897 VGND.n895 4.5005
R1532 VGND.n150 VGND.n149 4.5005
R1533 VGND.n925 VGND.n922 4.5005
R1534 VGND.n971 VGND.n970 4.5005
R1535 VGND.n930 VGND.n927 4.5005
R1536 VGND.n809 VGND.n169 4.5005
R1537 VGND.n817 VGND.n816 4.5005
R1538 VGND.n299 VGND.n298 4.5005
R1539 VGND.n287 VGND.n234 4.5005
R1540 VGND.n292 VGND.n291 4.5005
R1541 VGND.n1339 VGND.n1338 4.5005
R1542 VGND.n13 VGND.n12 4.5005
R1543 VGND.n4 VGND.n3 4.5005
R1544 VGND.n257 VGND.n30 4.5005
R1545 VGND.n1310 VGND.n1309 4.5005
R1546 VGND.n33 VGND.n32 4.5005
R1547 VGND.n991 VGND.n990 4.42603
R1548 VGND.n337 VGND.n336 4.38651
R1549 VGND.n378 VGND.n368 4.36875
R1550 VGND.n729 VGND.n312 4.36875
R1551 VGND.n729 VGND.n728 4.36875
R1552 VGND.n723 VGND.n313 4.36875
R1553 VGND.n508 VGND.n507 4.36875
R1554 VGND.n483 VGND.n472 4.36875
R1555 VGND.n536 VGND.n535 4.36875
R1556 VGND.n465 VGND.n464 4.36875
R1557 VGND.n946 VGND.n942 4.36875
R1558 VGND.n143 VGND.n142 4.36875
R1559 VGND.n953 VGND.n938 4.36875
R1560 VGND.n952 VGND.n951 4.36875
R1561 VGND.n968 VGND.n928 4.36875
R1562 VGND.n961 VGND.n937 4.36875
R1563 VGND.n364 VGND.n363 4.35795
R1564 VGND.n542 VGND.n541 4.35795
R1565 VGND.n554 VGND.n410 4.28986
R1566 VGND.n586 VGND.n585 4.28986
R1567 VGND.n989 VGND.n918 4.28986
R1568 VGND.n1217 VGND.n1206 4.14168
R1569 VGND.n195 VGND.n191 4.11798
R1570 VGND.n225 VGND.n195 4.11798
R1571 VGND.n688 VGND.n388 4.11798
R1572 VGND.n685 VGND.n388 4.11798
R1573 VGND.n601 VGND.n600 4.11798
R1574 VGND.n600 VGND.n599 4.11798
R1575 VGND.n1144 VGND.n123 4.11798
R1576 VGND.n1141 VGND.n123 4.11798
R1577 VGND.n1012 VGND.n1002 4.11798
R1578 VGND.n1013 VGND.n1012 4.11798
R1579 VGND.n585 VGND.n583 4.07323
R1580 VGND.n541 VGND.n447 4.04261
R1581 VGND.n1090 VGND.n1089 3.97459
R1582 VGND.n774 VGND.n773 3.96548
R1583 VGND.n981 VGND.n980 3.96548
R1584 VGND.n1060 VGND.n1059 3.93896
R1585 VGND.n1198 VGND.n1196 3.76521
R1586 VGND.n1061 VGND.n1060 3.75994
R1587 VGND.n693 VGND.n387 3.7575
R1588 VGND.n775 VGND.n774 3.7069
R1589 VGND.n981 VGND.n919 3.7069
R1590 VGND.n980 VGND.n979 3.7069
R1591 VGND.n773 VGND.n186 3.68605
R1592 VGND.n985 VGND.n984 3.59021
R1593 VGND.n861 VGND.n845 3.50735
R1594 VGND.n1176 VGND.n55 3.50735
R1595 VGND.n806 VGND.n805 3.48706
R1596 VGND.n350 VGND.n349 3.48706
R1597 VGND.n891 VGND.n890 3.48706
R1598 VGND.n900 VGND.n899 3.48706
R1599 VGND.n812 VGND.n811 3.48706
R1600 VGND.n425 VGND.n424 3.45831
R1601 VGND.n441 VGND.n438 3.44377
R1602 VGND.n912 VGND.n909 3.44377
R1603 VGND.n446 VGND.n445 3.44339
R1604 VGND.n290 VGND.n230 3.43925
R1605 VGND.n301 VGND.n300 3.43925
R1606 VGND.n1344 VGND.n1343 3.43925
R1607 VGND.n1341 VGND.n1340 3.43925
R1608 VGND.n1065 VGND.n1064 3.43925
R1609 VGND.n1069 VGND.n1068 3.43925
R1610 VGND.n1306 VGND.n1305 3.43925
R1611 VGND.n526 VGND.n525 3.43925
R1612 VGND.n530 VGND.n529 3.43925
R1613 VGND.n815 VGND.n814 3.43925
R1614 VGND.n1257 VGND.n1256 3.43925
R1615 VGND.n1214 VGND.n1213 3.43925
R1616 VGND.n1292 VGND.n36 3.43925
R1617 VGND.n1302 VGND.n1301 3.43925
R1618 VGND.n760 VGND.n759 3.43925
R1619 VGND.n757 VGND.n756 3.43925
R1620 VGND.n176 VGND.n172 3.43925
R1621 VGND.n668 VGND.n667 3.43925
R1622 VGND.n622 VGND.n621 3.43925
R1623 VGND.n703 VGND.n702 3.43925
R1624 VGND.n707 VGND.n706 3.43925
R1625 VGND.n736 VGND.n303 3.43925
R1626 VGND.n748 VGND.n747 3.43925
R1627 VGND.n354 VGND.n353 3.43925
R1628 VGND.n903 VGND.n902 3.43925
R1629 VGND.n156 VGND.n153 3.43925
R1630 VGND.n608 VGND.n402 3.43925
R1631 VGND.n618 VGND.n617 3.43925
R1632 VGND.n489 VGND.n488 3.43925
R1633 VGND.n479 VGND.n478 3.43925
R1634 VGND.n1098 VGND.n136 3.43925
R1635 VGND.n1108 VGND.n1107 3.43925
R1636 VGND.n258 VGND.n35 3.43925
R1637 VGND.n1159 VGND.n115 3.43925
R1638 VGND.n854 VGND.n114 3.43925
R1639 VGND.n112 VGND.n111 3.43925
R1640 VGND.n1165 VGND.n1164 3.43925
R1641 VGND.n233 VGND.n231 3.4105
R1642 VGND.n289 VGND.n288 3.4105
R1643 VGND.n9 VGND.n7 3.4105
R1644 VGND.n11 VGND.n5 3.4105
R1645 VGND.n1067 VGND.n1005 3.4105
R1646 VGND.n1066 VGND.n1006 3.4105
R1647 VGND.n528 VGND.n453 3.4105
R1648 VGND.n527 VGND.n454 3.4105
R1649 VGND.n810 VGND.n808 3.4105
R1650 VGND.n171 VGND.n170 3.4105
R1651 VGND.n1215 VGND.n1209 3.4105
R1652 VGND.n1259 VGND.n1258 3.4105
R1653 VGND.n40 VGND.n38 3.4105
R1654 VGND.n47 VGND.n46 3.4105
R1655 VGND.n752 VGND.n750 3.4105
R1656 VGND.n229 VGND.n193 3.4105
R1657 VGND.n804 VGND.n174 3.4105
R1658 VGND.n802 VGND.n801 3.4105
R1659 VGND.n401 VGND.n399 3.4105
R1660 VGND.n670 VGND.n669 3.4105
R1661 VGND.n705 VGND.n323 3.4105
R1662 VGND.n704 VGND.n324 3.4105
R1663 VGND.n307 VGND.n305 3.4105
R1664 VGND.n735 VGND.n734 3.4105
R1665 VGND.n351 VGND.n348 3.4105
R1666 VGND.n352 VGND.n346 3.4105
R1667 VGND.n898 VGND.n893 3.4105
R1668 VGND.n896 VGND.n151 3.4105
R1669 VGND.n889 VGND.n154 3.4105
R1670 VGND.n887 VGND.n886 3.4105
R1671 VGND.n431 VGND.n152 3.4105
R1672 VGND.n424 VGND.n152 3.4105
R1673 VGND.n432 VGND.n431 3.4105
R1674 VGND.n423 VGND.n422 3.4105
R1675 VGND.n430 VGND.n429 3.4105
R1676 VGND.n405 VGND.n403 3.4105
R1677 VGND.n607 VGND.n606 3.4105
R1678 VGND.n480 VGND.n475 3.4105
R1679 VGND.n491 VGND.n490 3.4105
R1680 VGND.n139 VGND.n137 3.4105
R1681 VGND.n1097 VGND.n1096 3.4105
R1682 VGND.n1124 VGND.n1114 3.4105
R1683 VGND.n1114 VGND.n1113 3.4105
R1684 VGND.n1124 VGND.n1123 3.4105
R1685 VGND.n1113 VGND.n1112 3.4105
R1686 VGND.n1110 VGND.n132 3.4105
R1687 VGND.n1126 VGND.n1125 3.4105
R1688 VGND.n852 VGND.n116 3.4105
R1689 VGND.n1158 VGND.n1157 3.4105
R1690 VGND.n68 VGND.n62 3.4105
R1691 VGND.n69 VGND.n64 3.4105
R1692 VGND.n932 VGND.n113 3.4105
R1693 VGND.n974 VGND.n113 3.4105
R1694 VGND.n933 VGND.n932 3.4105
R1695 VGND.n975 VGND.n974 3.4105
R1696 VGND.n973 VGND.n972 3.4105
R1697 VGND.n931 VGND.n924 3.4105
R1698 VGND.n34 VGND.n31 3.4105
R1699 VGND.n1308 VGND.n1307 3.4105
R1700 VGND.n699 VGND.n337 3.31239
R1701 VGND.n438 VGND.n437 3.21921
R1702 VGND.n909 VGND.n908 3.21921
R1703 VGND.n858 VGND.n857 3.2005
R1704 VGND.n1173 VGND.n1172 3.2005
R1705 VGND.n1296 VGND.n44 3.13241
R1706 VGND.n1120 VGND.n1119 3.13241
R1707 VGND.n830 VGND.n829 3.13241
R1708 VGND.n1091 VGND.n1090 3.05276
R1709 VGND.n1229 VGND.n1227 3.04861
R1710 VGND.n639 VGND.n637 3.04861
R1711 VGND.n581 VGND.n578 3.04861
R1712 VGND.n1034 VGND.n1032 3.04861
R1713 VGND.n583 VGND.n582 3.04861
R1714 VGND.n1018 VGND.n1011 3.04386
R1715 VGND.n693 VGND.n692 3.01483
R1716 VGND.n787 VGND.n786 2.99624
R1717 VGND.n557 VGND.n410 2.9514
R1718 VGND.n558 VGND.n557 2.9514
R1719 VGND.n562 VGND.n561 2.92131
R1720 VGND.n198 VGND.n197 2.77533
R1721 VGND.n786 VGND.n785 2.7239
R1722 VGND.n48 VGND.n44 2.7239
R1723 VGND.n1119 VGND.n1118 2.7239
R1724 VGND.n829 VGND.n165 2.7239
R1725 VGND.n847 VGND.n846 2.63064
R1726 VGND.n57 VGND.n56 2.63064
R1727 VGND.n769 VGND.n188 2.55412
R1728 VGND.n371 VGND.n369 2.33701
R1729 VGND.n372 VGND.n371 2.33701
R1730 VGND.n743 VGND.n742 2.33701
R1731 VGND.n317 VGND.n315 2.33701
R1732 VGND.n717 VGND.n317 2.33701
R1733 VGND.n715 VGND.n318 2.33701
R1734 VGND.n500 VGND.n470 2.33701
R1735 VGND.n497 VGND.n470 2.33701
R1736 VGND.n497 VGND.n496 2.33701
R1737 VGND.n496 VGND.n495 2.33701
R1738 VGND.n522 VGND.n521 2.33701
R1739 VGND.n521 VGND.n520 2.33701
R1740 VGND.n520 VGND.n519 2.33701
R1741 VGND.n519 VGND.n518 2.33701
R1742 VGND.n944 VGND.n141 2.33701
R1743 VGND.n1103 VGND.n141 2.33701
R1744 VGND.n936 VGND.n929 2.33701
R1745 VGND.n963 VGND.n936 2.33701
R1746 VGND.n805 VGND.n175 2.33488
R1747 VGND.n349 VGND.n344 2.33488
R1748 VGND.n427 VGND.n425 2.33488
R1749 VGND.n890 VGND.n155 2.33488
R1750 VGND.n899 VGND.n895 2.33488
R1751 VGND.n811 VGND.n169 2.33488
R1752 VGND.n768 VGND.n189 2.33067
R1753 VGND.n557 VGND.n556 2.25312
R1754 VGND.n363 VGND.n362 2.10893
R1755 VGND.n742 VGND.n741 2.03225
R1756 VGND.n319 VGND.n318 2.03225
R1757 VGND.n766 VGND.n765 1.91571
R1758 VGND.n990 VGND.n989 1.8388
R1759 VGND.n441 VGND.n440 1.72214
R1760 VGND.n912 VGND.n911 1.72214
R1761 VGND.n892 VGND.n153 1.69188
R1762 VGND.n892 VGND.n891 1.69188
R1763 VGND.n902 VGND.n901 1.69188
R1764 VGND.n901 VGND.n900 1.69188
R1765 VGND.n353 VGND.n173 1.69188
R1766 VGND.n350 VGND.n173 1.69188
R1767 VGND.n807 VGND.n172 1.69188
R1768 VGND.n807 VGND.n806 1.69188
R1769 VGND.n814 VGND.n813 1.69188
R1770 VGND.n813 VGND.n812 1.69188
R1771 VGND.n421 VGND.n152 1.69188
R1772 VGND.n1109 VGND.n136 1.69188
R1773 VGND.n1109 VGND.n1108 1.69188
R1774 VGND.n489 VGND.n135 1.69188
R1775 VGND.n479 VGND.n135 1.69188
R1776 VGND.n703 VGND.n37 1.69188
R1777 VGND.n706 VGND.n37 1.69188
R1778 VGND.n1303 VGND.n36 1.69188
R1779 VGND.n1303 VGND.n1302 1.69188
R1780 VGND.n1306 VGND.n1304 1.69188
R1781 VGND.n1304 VGND.n35 1.69188
R1782 VGND.n1114 VGND.n134 1.69188
R1783 VGND.n1163 VGND.n112 1.69188
R1784 VGND.n1164 VGND.n1163 1.69188
R1785 VGND.n1065 VGND.n63 1.69188
R1786 VGND.n1068 VGND.n63 1.69188
R1787 VGND.n619 VGND.n402 1.69188
R1788 VGND.n619 VGND.n618 1.69188
R1789 VGND.n668 VGND.n623 1.69188
R1790 VGND.n623 VGND.n622 1.69188
R1791 VGND.n1257 VGND.n6 1.69188
R1792 VGND.n1214 VGND.n6 1.69188
R1793 VGND.n1343 VGND.n1342 1.69188
R1794 VGND.n1342 VGND.n1341 1.69188
R1795 VGND.n1160 VGND.n114 1.69188
R1796 VGND.n1160 VGND.n1159 1.69188
R1797 VGND.n526 VGND.n304 1.69188
R1798 VGND.n529 VGND.n304 1.69188
R1799 VGND.n749 VGND.n303 1.69188
R1800 VGND.n749 VGND.n748 1.69188
R1801 VGND.n759 VGND.n758 1.69188
R1802 VGND.n758 VGND.n757 1.69188
R1803 VGND.n302 VGND.n230 1.69188
R1804 VGND.n302 VGND.n301 1.69188
R1805 VGND.n923 VGND.n113 1.69188
R1806 VGND.n918 VGND.n917 1.5365
R1807 VGND.n210 VGND.n204 1.50638
R1808 VGND.n440 VGND.n439 1.49758
R1809 VGND.n911 VGND.n910 1.49758
R1810 VGND.n485 VGND.n484 1.47352
R1811 VGND.n958 VGND.n957 1.46433
R1812 VGND.n957 VGND.n956 1.42881
R1813 VGND.n545 VGND.n445 1.3622
R1814 VGND.n776 VGND.n184 1.20723
R1815 VGND.n1357 VGND.n1356 1.18311
R1816 VGND.n265 VGND.n264 1.18311
R1817 VGND.n160 VGND.n159 1.18311
R1818 VGND.n87 VGND.n86 1.18311
R1819 VGND.n820 VGND.n819 1.18311
R1820 VGND.n857 VGND.n846 1.14023
R1821 VGND.n1172 VGND.n56 1.14023
R1822 VGND.n1218 VGND.n1217 1.12991
R1823 VGND.n585 VGND.n584 0.952566
R1824 VGND.n583 VGND.n580 0.899674
R1825 VGND.n643 VGND.n642 0.835283
R1826 VGND.n1038 VGND.n1037 0.835283
R1827 VGND.n858 VGND.n845 0.833377
R1828 VGND.n1173 VGND.n55 0.833377
R1829 VGND.n766 VGND.n189 0.830425
R1830 VGND.n1053 VGND.n1052 0.753441
R1831 VGND.n692 VGND.n691 0.743162
R1832 VGND.n410 VGND.n409 0.69032
R1833 VGND.n559 VGND.n558 0.69032
R1834 VGND.n769 VGND.n768 0.606984
R1835 VGND.n220 VGND.n198 0.537563
R1836 VGND.n680 VGND.n390 0.537563
R1837 VGND.n336 VGND.n335 0.537563
R1838 VGND.n330 VGND.n329 0.537563
R1839 VGND.n594 VGND.n593 0.537563
R1840 VGND.n848 VGND.n120 0.537563
R1841 VGND.n1136 VGND.n125 0.537563
R1842 VGND.n1081 VGND.n997 0.537563
R1843 VGND.n1000 VGND.n998 0.537563
R1844 VGND.n1059 VGND.n1058 0.537563
R1845 VGND.n1085 VGND.n1084 0.537563
R1846 VGND.n1083 VGND.n1082 0.537563
R1847 VGND.n862 VGND.n861 0.526527
R1848 VGND.n1177 VGND.n1176 0.526527
R1849 VGND.n1360 VGND.n1359 0.417891
R1850 VGND.n268 VGND.n267 0.417891
R1851 VGND.n264 VGND.n263 0.417891
R1852 VGND.n647 VGND.n634 0.417891
R1853 VGND.n641 VGND.n640 0.417891
R1854 VGND.n880 VGND.n879 0.417891
R1855 VGND.n90 VGND.n89 0.417891
R1856 VGND.n1042 VGND.n1029 0.417891
R1857 VGND.n1036 VGND.n1035 0.417891
R1858 VGND.n821 VGND.n167 0.417891
R1859 VGND.n792 VGND.n177 0.409011
R1860 VGND.n785 VGND.n784 0.409011
R1861 VGND.n205 VGND.n43 0.409011
R1862 VGND.n1289 VGND.n48 0.409011
R1863 VGND.n361 VGND.n360 0.409011
R1864 VGND.n553 VGND.n552 0.409011
R1865 VGND.n591 VGND.n573 0.409011
R1866 VGND.n869 VGND.n868 0.409011
R1867 VGND.n1130 VGND.n129 0.409011
R1868 VGND.n1118 VGND.n49 0.409011
R1869 VGND.n1184 VGND.n1183 0.409011
R1870 VGND.n827 VGND.n826 0.409011
R1871 VGND.n833 VGND.n165 0.409011
R1872 VGND.n188 VGND.n186 0.383542
R1873 VGND.n651 VGND.n650 0.376971
R1874 VGND.n657 VGND.n655 0.376971
R1875 VGND.n1046 VGND.n1045 0.376971
R1876 VGND.n642 VGND.n641 0.348326
R1877 VGND.n1037 VGND.n1036 0.348326
R1878 VGND.n179 VGND.n177 0.340926
R1879 VGND.n368 VGND.n339 0.305262
R1880 VGND.n741 VGND.n740 0.305262
R1881 VGND.n312 VGND.n310 0.305262
R1882 VGND.n728 VGND.n727 0.305262
R1883 VGND.n726 VGND.n313 0.305262
R1884 VGND.n712 VGND.n319 0.305262
R1885 VGND.n509 VGND.n508 0.305262
R1886 VGND.n485 VGND.n483 0.305262
R1887 VGND.n537 VGND.n536 0.305262
R1888 VGND.n514 VGND.n465 0.305262
R1889 VGND.n942 VGND.n940 0.305262
R1890 VGND.n1091 VGND.n143 0.305262
R1891 VGND.n956 VGND.n938 0.305262
R1892 VGND.n951 VGND.n950 0.305262
R1893 VGND.n928 VGND.n921 0.305262
R1894 VGND.n958 VGND.n937 0.305262
R1895 VGND.n689 VGND.n688 0.269031
R1896 VGND.n593 VGND.n592 0.269031
R1897 VGND.n849 VGND.n847 0.263514
R1898 VGND.n1169 VGND.n57 0.263514
R1899 VGND.n387 VGND.n385 0.262616
R1900 VGND.n691 VGND.n690 0.262616
R1901 VGND.n776 VGND.n775 0.259086
R1902 VGND.n984 VGND.n919 0.259086
R1903 VGND.n979 VGND.n978 0.259086
R1904 VGND.n1161 VGND 0.241669
R1905 VGND VGND.n1162 0.241669
R1906 VGND.n582 VGND.n574 0.239726
R1907 VGND.n556 VGND 0.238178
R1908 VGND.n437 VGND.n436 0.225061
R1909 VGND.n439 VGND.n414 0.225061
R1910 VGND.n908 VGND.n907 0.225061
R1911 VGND.n910 VGND.n144 0.225061
R1912 VGND.n1162 VGND.n1161 0.2167
R1913 VGND.n556 VGND 0.199635
R1914 VGND.n765 VGND.n764 0.192021
R1915 VGND.n602 VGND.n569 0.179521
R1916 VGND.n1227 VGND 0.179485
R1917 VGND.n637 VGND 0.179485
R1918 VGND VGND.n581 0.179485
R1919 VGND.n1032 VGND 0.179485
R1920 VGND.n813 VGND.n807 0.1603
R1921 VGND.n807 VGND.n173 0.1603
R1922 VGND.n173 VGND.n152 0.1603
R1923 VGND.n901 VGND.n152 0.1603
R1924 VGND.n901 VGND.n892 0.1603
R1925 VGND.n1304 VGND.n1303 0.1603
R1926 VGND.n1303 VGND.n37 0.1603
R1927 VGND.n135 VGND.n37 0.1603
R1928 VGND.n1109 VGND.n135 0.1603
R1929 VGND.n1114 VGND.n1109 0.1603
R1930 VGND.n1342 VGND.n6 0.1603
R1931 VGND.n623 VGND.n6 0.1603
R1932 VGND.n623 VGND.n619 0.1603
R1933 VGND.n619 VGND.n63 0.1603
R1934 VGND.n1163 VGND.n63 0.1603
R1935 VGND.n758 VGND.n302 0.1603
R1936 VGND.n758 VGND.n749 0.1603
R1937 VGND.n749 VGND.n304 0.1603
R1938 VGND.n304 VGND.n113 0.1603
R1939 VGND.n1160 VGND.n113 0.1603
R1940 VGND.n1227 VGND 0.14207
R1941 VGND.n637 VGND 0.14207
R1942 VGND.n581 VGND 0.14207
R1943 VGND.n1032 VGND 0.14207
R1944 VGND.n582 VGND 0.141725
R1945 VGND.n788 VGND.n787 0.13667
R1946 VGND.n797 VGND 0.120408
R1947 VGND.n343 VGND 0.120408
R1948 VGND VGND.n434 0.120408
R1949 VGND VGND.n905 0.120408
R1950 VGND.n366 VGND 0.120408
R1951 VGND.n564 VGND 0.120408
R1952 VGND VGND.n987 0.120408
R1953 VGND.n791 VGND.n790 0.120292
R1954 VGND.n790 VGND.n178 0.120292
R1955 VGND.n783 VGND.n178 0.120292
R1956 VGND.n777 VGND.n185 0.120292
R1957 VGND.n772 VGND.n185 0.120292
R1958 VGND.n772 VGND.n771 0.120292
R1959 VGND.n771 VGND.n770 0.120292
R1960 VGND.n227 VGND.n226 0.120292
R1961 VGND.n226 VGND.n194 0.120292
R1962 VGND.n222 VGND.n194 0.120292
R1963 VGND.n222 VGND.n221 0.120292
R1964 VGND.n217 VGND.n216 0.120292
R1965 VGND.n213 VGND.n212 0.120292
R1966 VGND.n212 VGND.n211 0.120292
R1967 VGND.n211 VGND.n202 0.120292
R1968 VGND.n1280 VGND.n1279 0.120292
R1969 VGND.n1269 VGND.n1268 0.120292
R1970 VGND.n1268 VGND.n1205 0.120292
R1971 VGND.n1250 VGND.n1249 0.120292
R1972 VGND.n1249 VGND.n1248 0.120292
R1973 VGND.n1248 VGND.n1221 0.120292
R1974 VGND.n1242 VGND.n1221 0.120292
R1975 VGND.n1235 VGND.n1234 0.120292
R1976 VGND.n1234 VGND.n1233 0.120292
R1977 VGND.n1233 VGND.n1225 0.120292
R1978 VGND.n365 VGND.n341 0.120292
R1979 VGND.n380 VGND.n379 0.120292
R1980 VGND.n379 VGND.n367 0.120292
R1981 VGND.n375 VGND.n367 0.120292
R1982 VGND.n375 VGND.n374 0.120292
R1983 VGND.n374 VGND.n373 0.120292
R1984 VGND.n373 VGND.n370 0.120292
R1985 VGND.n731 VGND.n730 0.120292
R1986 VGND.n730 VGND.n311 0.120292
R1987 VGND.n725 VGND.n724 0.120292
R1988 VGND.n724 VGND.n314 0.120292
R1989 VGND.n720 VGND.n314 0.120292
R1990 VGND.n720 VGND.n719 0.120292
R1991 VGND.n719 VGND.n718 0.120292
R1992 VGND.n718 VGND.n316 0.120292
R1993 VGND.n714 VGND.n316 0.120292
R1994 VGND.n714 VGND.n713 0.120292
R1995 VGND.n710 VGND.n709 0.120292
R1996 VGND.n700 VGND.n327 0.120292
R1997 VGND.n695 VGND.n694 0.120292
R1998 VGND.n694 VGND.n386 0.120292
R1999 VGND.n686 VGND.n389 0.120292
R2000 VGND.n682 VGND.n389 0.120292
R2001 VGND.n682 VGND.n681 0.120292
R2002 VGND.n678 VGND.n677 0.120292
R2003 VGND.n665 VGND.n625 0.120292
R2004 VGND.n661 VGND.n625 0.120292
R2005 VGND.n659 VGND.n628 0.120292
R2006 VGND.n652 VGND.n631 0.120292
R2007 VGND.n646 VGND.n645 0.120292
R2008 VGND.n645 VGND.n635 0.120292
R2009 VGND.n435 VGND.n415 0.120292
R2010 VGND.n442 VGND.n415 0.120292
R2011 VGND.n443 VGND.n442 0.120292
R2012 VGND.n544 VGND.n543 0.120292
R2013 VGND.n538 VGND.n449 0.120292
R2014 VGND.n533 VGND.n449 0.120292
R2015 VGND.n533 VGND.n532 0.120292
R2016 VGND.n523 VGND.n457 0.120292
R2017 VGND.n517 VGND.n457 0.120292
R2018 VGND.n517 VGND.n516 0.120292
R2019 VGND.n516 VGND.n515 0.120292
R2020 VGND.n510 VGND.n467 0.120292
R2021 VGND.n505 VGND.n467 0.120292
R2022 VGND.n505 VGND.n504 0.120292
R2023 VGND.n504 VGND.n503 0.120292
R2024 VGND.n503 VGND.n469 0.120292
R2025 VGND.n499 VGND.n469 0.120292
R2026 VGND.n499 VGND.n498 0.120292
R2027 VGND.n603 VGND.n570 0.120292
R2028 VGND.n598 VGND.n570 0.120292
R2029 VGND.n598 VGND.n597 0.120292
R2030 VGND.n597 VGND.n596 0.120292
R2031 VGND.n596 VGND.n572 0.120292
R2032 VGND.n589 VGND.n574 0.120292
R2033 VGND.n882 VGND.n157 0.120292
R2034 VGND.n876 VGND.n875 0.120292
R2035 VGND.n870 VGND.n842 0.120292
R2036 VGND.n865 VGND.n842 0.120292
R2037 VGND.n865 VGND.n864 0.120292
R2038 VGND.n864 VGND.n863 0.120292
R2039 VGND.n863 VGND.n844 0.120292
R2040 VGND.n856 VGND.n844 0.120292
R2041 VGND.n1153 VGND.n119 0.120292
R2042 VGND.n1149 VGND.n119 0.120292
R2043 VGND.n1149 VGND.n1148 0.120292
R2044 VGND.n1148 VGND.n1147 0.120292
R2045 VGND.n1147 VGND.n122 0.120292
R2046 VGND.n1143 VGND.n122 0.120292
R2047 VGND.n1143 VGND.n1142 0.120292
R2048 VGND.n1142 VGND.n124 0.120292
R2049 VGND.n1138 VGND.n124 0.120292
R2050 VGND.n1138 VGND.n1137 0.120292
R2051 VGND.n1133 VGND.n1132 0.120292
R2052 VGND.n1121 VGND.n1116 0.120292
R2053 VGND.n1187 VGND.n1186 0.120292
R2054 VGND.n1185 VGND.n52 0.120292
R2055 VGND.n1180 VGND.n52 0.120292
R2056 VGND.n1180 VGND.n1179 0.120292
R2057 VGND.n1179 VGND.n1178 0.120292
R2058 VGND.n1178 VGND.n54 0.120292
R2059 VGND.n1171 VGND.n54 0.120292
R2060 VGND.n1171 VGND.n1170 0.120292
R2061 VGND.n109 VGND.n66 0.120292
R2062 VGND.n76 VGND.n66 0.120292
R2063 VGND.n104 VGND.n76 0.120292
R2064 VGND.n104 VGND.n103 0.120292
R2065 VGND.n103 VGND.n102 0.120292
R2066 VGND.n98 VGND.n97 0.120292
R2067 VGND.n97 VGND.n81 0.120292
R2068 VGND.n93 VGND.n81 0.120292
R2069 VGND.n93 VGND.n92 0.120292
R2070 VGND.n91 VGND.n84 0.120292
R2071 VGND.n85 VGND.n84 0.120292
R2072 VGND.n906 VGND.n145 0.120292
R2073 VGND.n913 VGND.n145 0.120292
R2074 VGND.n914 VGND.n913 0.120292
R2075 VGND.n983 VGND.n982 0.120292
R2076 VGND.n982 VGND.n920 0.120292
R2077 VGND.n977 VGND.n920 0.120292
R2078 VGND.n966 VGND.n965 0.120292
R2079 VGND.n965 VGND.n964 0.120292
R2080 VGND.n964 VGND.n935 0.120292
R2081 VGND.n960 VGND.n935 0.120292
R2082 VGND.n960 VGND.n959 0.120292
R2083 VGND.n955 VGND.n954 0.120292
R2084 VGND.n954 VGND.n939 0.120292
R2085 VGND.n949 VGND.n939 0.120292
R2086 VGND.n948 VGND.n947 0.120292
R2087 VGND.n947 VGND.n941 0.120292
R2088 VGND.n943 VGND.n941 0.120292
R2089 VGND.n1093 VGND.n1092 0.120292
R2090 VGND.n1086 VGND.n995 0.120292
R2091 VGND.n1080 VGND 0.120292
R2092 VGND.n1076 VGND.n1075 0.120292
R2093 VGND.n1075 VGND.n999 0.120292
R2094 VGND VGND.n999 0.120292
R2095 VGND.n1062 VGND.n1009 0.120292
R2096 VGND.n1055 VGND.n1054 0.120292
R2097 VGND.n1054 VGND.n1021 0.120292
R2098 VGND.n1047 VGND.n1026 0.120292
R2099 VGND.n1041 VGND.n1040 0.120292
R2100 VGND.n1040 VGND.n1030 0.120292
R2101 VGND.n824 VGND.n823 0.120292
R2102 VGND.n825 VGND.n166 0.120292
R2103 VGND.n831 VGND.n166 0.120292
R2104 VGND.n832 VGND.n831 0.120292
R2105 VGND.n241 VGND.n240 0.120292
R2106 VGND.n241 VGND.n238 0.120292
R2107 VGND.n245 VGND.n238 0.120292
R2108 VGND.n246 VGND.n245 0.120292
R2109 VGND.n247 VGND.n246 0.120292
R2110 VGND.n285 VGND.n284 0.120292
R2111 VGND.n284 VGND.n251 0.120292
R2112 VGND.n279 VGND.n278 0.120292
R2113 VGND.n278 VGND.n277 0.120292
R2114 VGND.n277 VGND.n253 0.120292
R2115 VGND.n271 VGND.n253 0.120292
R2116 VGND.n271 VGND.n270 0.120292
R2117 VGND.n269 VGND.n255 0.120292
R2118 VGND.n262 VGND.n255 0.120292
R2119 VGND.n1316 VGND.n1315 0.120292
R2120 VGND.n1322 VGND.n1321 0.120292
R2121 VGND.n1327 VGND.n1326 0.120292
R2122 VGND.n1327 VGND.n17 0.120292
R2123 VGND.n1331 VGND.n17 0.120292
R2124 VGND.n1332 VGND.n1331 0.120292
R2125 VGND.n1346 VGND.n0 0.120292
R2126 VGND.n1375 VGND.n1374 0.120292
R2127 VGND.n1369 VGND.n1368 0.120292
R2128 VGND.n1368 VGND.n1352 0.120292
R2129 VGND.n1363 VGND.n1352 0.120292
R2130 VGND.n1363 VGND.n1362 0.120292
R2131 VGND.n1361 VGND.n1354 0.120292
R2132 VGND.n1355 VGND.n1354 0.120292
R2133 VGND.n1235 VGND 0.0994583
R2134 VGND.n218 VGND 0.0981562
R2135 VGND VGND.n1280 0.0981562
R2136 VGND VGND.n1269 0.0981562
R2137 VGND.n1250 VGND 0.0981562
R2138 VGND.n725 VGND 0.0981562
R2139 VGND.n710 VGND 0.0981562
R2140 VGND.n678 VGND 0.0981562
R2141 VGND VGND.n652 0.0981562
R2142 VGND.n511 VGND 0.0981562
R2143 VGND VGND.n510 0.0981562
R2144 VGND VGND.n482 0.0981562
R2145 VGND.n550 VGND 0.0981562
R2146 VGND.n566 VGND 0.0981562
R2147 VGND VGND.n589 0.0981562
R2148 VGND.n1134 VGND 0.0981562
R2149 VGND VGND.n98 0.0981562
R2150 VGND.n955 VGND 0.0981562
R2151 VGND VGND.n948 0.0981562
R2152 VGND.n1088 VGND 0.0981562
R2153 VGND.n1080 VGND 0.0981562
R2154 VGND.n1056 VGND 0.0981562
R2155 VGND VGND.n1047 0.0981562
R2156 VGND VGND.n260 0.0981562
R2157 VGND.n1321 VGND 0.0981562
R2158 VGND.n1326 VGND 0.0981562
R2159 VGND VGND.n14 0.0981562
R2160 VGND.n1375 VGND 0.0981562
R2161 VGND VGND.n1369 0.0981562
R2162 VGND VGND.n686 0.0968542
R2163 VGND VGND.n876 0.0955521
R2164 VGND VGND.n1133 0.0955521
R2165 VGND.n300 VGND.n299 0.0950946
R2166 VGND.n291 VGND.n290 0.0950946
R2167 VGND.n1340 VGND.n1339 0.0950946
R2168 VGND.n1344 VGND.n4 0.0950946
R2169 VGND.n1069 VGND.n1004 0.0950946
R2170 VGND.n1064 VGND.n1007 0.0950946
R2171 VGND.n530 VGND.n452 0.0950946
R2172 VGND.n525 VGND.n455 0.0950946
R2173 VGND.n816 VGND.n815 0.0950946
R2174 VGND.n1213 VGND.n1212 0.0950946
R2175 VGND.n1256 VGND.n1210 0.0950946
R2176 VGND.n1301 VGND.n1300 0.0950946
R2177 VGND.n1293 VGND.n1292 0.0950946
R2178 VGND.n756 VGND.n755 0.0950946
R2179 VGND.n761 VGND.n760 0.0950946
R2180 VGND.n800 VGND.n176 0.0950946
R2181 VGND.n621 VGND.n620 0.0950946
R2182 VGND.n667 VGND.n400 0.0950946
R2183 VGND.n707 VGND.n322 0.0950946
R2184 VGND.n702 VGND.n325 0.0950946
R2185 VGND.n747 VGND.n746 0.0950946
R2186 VGND.n737 VGND.n736 0.0950946
R2187 VGND.n355 VGND.n354 0.0950946
R2188 VGND.n903 VGND.n150 0.0950946
R2189 VGND.n885 VGND.n156 0.0950946
R2190 VGND.n432 VGND.n420 0.0950946
R2191 VGND.n617 VGND.n616 0.0950946
R2192 VGND.n609 VGND.n608 0.0950946
R2193 VGND.n478 VGND.n477 0.0950946
R2194 VGND.n488 VGND.n476 0.0950946
R2195 VGND.n1107 VGND.n1106 0.0950946
R2196 VGND.n1099 VGND.n1098 0.0950946
R2197 VGND.n1112 VGND.n1111 0.0950946
R2198 VGND.n1123 VGND.n133 0.0950946
R2199 VGND.n854 VGND.n853 0.0950946
R2200 VGND.n1156 VGND.n115 0.0950946
R2201 VGND.n1165 VGND.n61 0.0950946
R2202 VGND.n111 VGND.n65 0.0950946
R2203 VGND.n975 VGND.n922 0.0950946
R2204 VGND.n933 VGND.n930 0.0950946
R2205 VGND.n1305 VGND.n33 0.0950946
R2206 VGND.n811 VGND.n810 0.0878527
R2207 VGND.n805 VGND.n804 0.0878527
R2208 VGND.n349 VGND.n348 0.0878527
R2209 VGND.n899 VGND.n898 0.0878527
R2210 VGND.n890 VGND.n889 0.0878527
R2211 VGND.n425 VGND.n422 0.0878527
R2212 VGND.n799 VGND.n798 0.0838333
R2213 VGND.n754 VGND.n187 0.0838333
R2214 VGND.n1299 VGND.n39 0.0838333
R2215 VGND.n1211 VGND.n1207 0.0838333
R2216 VGND.n356 VGND.n345 0.0838333
R2217 VGND.n745 VGND.n306 0.0838333
R2218 VGND.n738 VGND.n732 0.0838333
R2219 VGND.n708 VGND.n321 0.0838333
R2220 VGND.n701 VGND.n326 0.0838333
R2221 VGND.n666 VGND.n624 0.0838333
R2222 VGND.n433 VGND.n419 0.0838333
R2223 VGND.n531 VGND.n451 0.0838333
R2224 VGND.n524 VGND.n456 0.0838333
R2225 VGND.n473 VGND.n471 0.0838333
R2226 VGND.n487 VGND.n481 0.0838333
R2227 VGND.n615 VGND.n404 0.0838333
R2228 VGND.n610 VGND.n604 0.0838333
R2229 VGND.n884 VGND.n883 0.0838333
R2230 VGND.n855 VGND.n851 0.0838333
R2231 VGND.n1155 VGND.n1154 0.0838333
R2232 VGND.n1122 VGND.n1115 0.0838333
R2233 VGND.n1166 VGND.n60 0.0838333
R2234 VGND.n904 VGND.n149 0.0838333
R2235 VGND.n934 VGND.n927 0.0838333
R2236 VGND.n1105 VGND.n138 0.0838333
R2237 VGND.n1100 VGND.n1094 0.0838333
R2238 VGND.n1070 VGND.n1003 0.0838333
R2239 VGND.n1063 VGND.n1008 0.0838333
R2240 VGND.n817 VGND.n168 0.0838333
R2241 VGND.n298 VGND.n232 0.0838333
R2242 VGND.n292 VGND.n286 0.0838333
R2243 VGND.n259 VGND.n30 0.0838333
R2244 VGND.n32 VGND.n25 0.0838333
R2245 VGND.n1338 VGND.n8 0.0838333
R2246 VGND.n1345 VGND.n3 0.0838333
R2247 VGND VGND.n366 0.082648
R2248 VGND VGND.n564 0.082648
R2249 VGND.n987 VGND 0.082648
R2250 VGND.n798 VGND.n797 0.0735334
R2251 VGND.n345 VGND.n343 0.0735334
R2252 VGND.n434 VGND.n433 0.0735334
R2253 VGND.n905 VGND.n904 0.0735334
R2254 VGND.n648 VGND.n647 0.0700652
R2255 VGND.n1043 VGND.n1042 0.0700652
R2256 VGND.n588 VGND.n587 0.0685851
R2257 VGND.n287 VGND.n233 0.0680676
R2258 VGND.n289 VGND.n287 0.0680676
R2259 VGND.n12 VGND.n9 0.0680676
R2260 VGND.n12 VGND.n11 0.0680676
R2261 VGND.n1015 VGND.n1005 0.0680676
R2262 VGND.n1015 VGND.n1006 0.0680676
R2263 VGND.n460 VGND.n453 0.0680676
R2264 VGND.n460 VGND.n454 0.0680676
R2265 VGND.n810 VGND.n809 0.0680676
R2266 VGND.n809 VGND.n170 0.0680676
R2267 VGND.n1260 VGND.n1209 0.0680676
R2268 VGND.n1260 VGND.n1259 0.0680676
R2269 VGND.n45 VGND.n40 0.0680676
R2270 VGND.n47 VGND.n45 0.0680676
R2271 VGND.n752 VGND.n751 0.0680676
R2272 VGND.n751 VGND.n193 0.0680676
R2273 VGND.n804 VGND.n803 0.0680676
R2274 VGND.n803 VGND.n802 0.0680676
R2275 VGND.n671 VGND.n399 0.0680676
R2276 VGND.n671 VGND.n670 0.0680676
R2277 VGND.n332 VGND.n323 0.0680676
R2278 VGND.n332 VGND.n324 0.0680676
R2279 VGND.n733 VGND.n307 0.0680676
R2280 VGND.n735 VGND.n733 0.0680676
R2281 VGND.n348 VGND.n347 0.0680676
R2282 VGND.n347 VGND.n346 0.0680676
R2283 VGND.n898 VGND.n897 0.0680676
R2284 VGND.n897 VGND.n896 0.0680676
R2285 VGND.n889 VGND.n888 0.0680676
R2286 VGND.n888 VGND.n887 0.0680676
R2287 VGND.n428 VGND.n422 0.0680676
R2288 VGND.n429 VGND.n428 0.0680676
R2289 VGND.n605 VGND.n405 0.0680676
R2290 VGND.n607 VGND.n605 0.0680676
R2291 VGND.n492 VGND.n475 0.0680676
R2292 VGND.n492 VGND.n491 0.0680676
R2293 VGND.n1095 VGND.n139 0.0680676
R2294 VGND.n1097 VGND.n1095 0.0680676
R2295 VGND.n1127 VGND.n132 0.0680676
R2296 VGND.n1127 VGND.n1126 0.0680676
R2297 VGND.n852 VGND.n117 0.0680676
R2298 VGND.n1157 VGND.n117 0.0680676
R2299 VGND.n70 VGND.n68 0.0680676
R2300 VGND.n70 VGND.n69 0.0680676
R2301 VGND.n972 VGND.n971 0.0680676
R2302 VGND.n971 VGND.n924 0.0680676
R2303 VGND.n258 VGND 0.0680676
R2304 VGND.n1309 VGND.n31 0.0680676
R2305 VGND.n1309 VGND.n1308 0.0680676
R2306 VGND.n795 VGND.n175 0.0603958
R2307 VGND.n791 VGND 0.0603958
R2308 VGND VGND.n782 0.0603958
R2309 VGND VGND.n781 0.0603958
R2310 VGND.n778 VGND 0.0603958
R2311 VGND VGND.n777 0.0603958
R2312 VGND.n753 VGND.n192 0.0603958
R2313 VGND.n763 VGND.n192 0.0603958
R2314 VGND VGND.n217 0.0603958
R2315 VGND.n216 VGND 0.0603958
R2316 VGND.n213 VGND 0.0603958
R2317 VGND.n207 VGND 0.0603958
R2318 VGND VGND.n206 0.0603958
R2319 VGND.n1298 VGND.n41 0.0603958
R2320 VGND.n1295 VGND.n41 0.0603958
R2321 VGND.n1287 VGND 0.0603958
R2322 VGND VGND.n1286 0.0603958
R2323 VGND VGND.n1285 0.0603958
R2324 VGND.n1281 VGND 0.0603958
R2325 VGND.n1279 VGND 0.0603958
R2326 VGND.n1276 VGND 0.0603958
R2327 VGND VGND.n1275 0.0603958
R2328 VGND VGND.n1274 0.0603958
R2329 VGND.n1274 VGND 0.0603958
R2330 VGND.n1270 VGND 0.0603958
R2331 VGND.n1262 VGND.n1261 0.0603958
R2332 VGND.n1261 VGND.n1208 0.0603958
R2333 VGND.n1242 VGND 0.0603958
R2334 VGND VGND.n1241 0.0603958
R2335 VGND VGND.n1240 0.0603958
R2336 VGND VGND.n1225 0.0603958
R2337 VGND.n357 VGND.n344 0.0603958
R2338 VGND VGND.n341 0.0603958
R2339 VGND.n381 VGND 0.0603958
R2340 VGND VGND.n380 0.0603958
R2341 VGND.n744 VGND.n308 0.0603958
R2342 VGND.n739 VGND.n308 0.0603958
R2343 VGND.n334 VGND.n333 0.0603958
R2344 VGND.n696 VGND 0.0603958
R2345 VGND VGND.n695 0.0603958
R2346 VGND.n687 VGND 0.0603958
R2347 VGND.n677 VGND 0.0603958
R2348 VGND VGND.n676 0.0603958
R2349 VGND.n673 VGND.n672 0.0603958
R2350 VGND.n672 VGND.n398 0.0603958
R2351 VGND VGND.n660 0.0603958
R2352 VGND.n660 VGND 0.0603958
R2353 VGND VGND.n659 0.0603958
R2354 VGND.n653 VGND 0.0603958
R2355 VGND.n646 VGND 0.0603958
R2356 VGND.n427 VGND.n426 0.0603958
R2357 VGND.n435 VGND 0.0603958
R2358 VGND.n444 VGND 0.0603958
R2359 VGND.n544 VGND 0.0603958
R2360 VGND.n539 VGND 0.0603958
R2361 VGND VGND.n538 0.0603958
R2362 VGND.n461 VGND.n459 0.0603958
R2363 VGND.n462 VGND.n461 0.0603958
R2364 VGND.n494 VGND.n493 0.0603958
R2365 VGND.n493 VGND.n474 0.0603958
R2366 VGND.n551 VGND 0.0603958
R2367 VGND.n555 VGND 0.0603958
R2368 VGND.n565 VGND 0.0603958
R2369 VGND.n614 VGND 0.0603958
R2370 VGND.n611 VGND 0.0603958
R2371 VGND.n590 VGND 0.0603958
R2372 VGND.n158 VGND.n155 0.0603958
R2373 VGND VGND.n157 0.0603958
R2374 VGND.n877 VGND 0.0603958
R2375 VGND.n875 VGND 0.0603958
R2376 VGND.n872 VGND 0.0603958
R2377 VGND VGND.n871 0.0603958
R2378 VGND VGND.n870 0.0603958
R2379 VGND VGND.n118 0.0603958
R2380 VGND.n1129 VGND.n1128 0.0603958
R2381 VGND.n1128 VGND.n131 0.0603958
R2382 VGND VGND.n50 0.0603958
R2383 VGND.n1187 VGND 0.0603958
R2384 VGND VGND.n1185 0.0603958
R2385 VGND.n1167 VGND 0.0603958
R2386 VGND.n71 VGND.n67 0.0603958
R2387 VGND.n73 VGND.n71 0.0603958
R2388 VGND.n99 VGND 0.0603958
R2389 VGND.n92 VGND 0.0603958
R2390 VGND VGND.n91 0.0603958
R2391 VGND.n895 VGND.n894 0.0603958
R2392 VGND.n906 VGND 0.0603958
R2393 VGND.n915 VGND 0.0603958
R2394 VGND.n988 VGND 0.0603958
R2395 VGND.n983 VGND 0.0603958
R2396 VGND.n970 VGND.n926 0.0603958
R2397 VGND.n970 VGND.n969 0.0603958
R2398 VGND.n1104 VGND.n140 0.0603958
R2399 VGND.n1101 VGND.n140 0.0603958
R2400 VGND VGND.n1087 0.0603958
R2401 VGND VGND.n1086 0.0603958
R2402 VGND.n1077 VGND 0.0603958
R2403 VGND VGND.n1076 0.0603958
R2404 VGND VGND.n1071 0.0603958
R2405 VGND.n1016 VGND.n1014 0.0603958
R2406 VGND.n1017 VGND.n1016 0.0603958
R2407 VGND VGND.n1055 0.0603958
R2408 VGND.n1048 VGND 0.0603958
R2409 VGND.n1041 VGND 0.0603958
R2410 VGND.n818 VGND.n169 0.0603958
R2411 VGND VGND.n824 0.0603958
R2412 VGND.n825 VGND 0.0603958
R2413 VGND VGND.n164 0.0603958
R2414 VGND.n240 VGND 0.0603958
R2415 VGND VGND.n235 0.0603958
R2416 VGND.n297 VGND.n234 0.0603958
R2417 VGND.n293 VGND.n234 0.0603958
R2418 VGND.n279 VGND 0.0603958
R2419 VGND VGND.n269 0.0603958
R2420 VGND VGND.n261 0.0603958
R2421 VGND.n1311 VGND.n1310 0.0603958
R2422 VGND.n1310 VGND.n26 0.0603958
R2423 VGND VGND.n1316 0.0603958
R2424 VGND.n1317 VGND 0.0603958
R2425 VGND.n1320 VGND 0.0603958
R2426 VGND.n1322 VGND 0.0603958
R2427 VGND.n1325 VGND 0.0603958
R2428 VGND VGND.n1332 0.0603958
R2429 VGND.n1333 VGND 0.0603958
R2430 VGND.n1337 VGND.n13 0.0603958
R2431 VGND.n13 VGND.n10 0.0603958
R2432 VGND VGND.n0 0.0603958
R2433 VGND VGND.n1379 0.0603958
R2434 VGND.n1374 VGND 0.0603958
R2435 VGND VGND.n1373 0.0603958
R2436 VGND.n1370 VGND 0.0603958
R2437 VGND.n1362 VGND 0.0603958
R2438 VGND VGND.n1361 0.0603958
R2439 VGND.n288 VGND.n231 0.0574697
R2440 VGND.n7 VGND.n5 0.0574697
R2441 VGND.n1067 VGND.n1066 0.0574697
R2442 VGND.n1307 VGND.n34 0.0574697
R2443 VGND.n528 VGND.n527 0.0574697
R2444 VGND.n808 VGND.n171 0.0574697
R2445 VGND.n1258 VGND.n1215 0.0574697
R2446 VGND.n46 VGND.n38 0.0574697
R2447 VGND.n750 VGND.n229 0.0574697
R2448 VGND.n801 VGND.n174 0.0574697
R2449 VGND.n669 VGND.n401 0.0574697
R2450 VGND.n705 VGND.n704 0.0574697
R2451 VGND.n734 VGND.n305 0.0574697
R2452 VGND.n352 VGND.n351 0.0574697
R2453 VGND.n893 VGND.n151 0.0574697
R2454 VGND.n886 VGND.n154 0.0574697
R2455 VGND.n424 VGND.n423 0.0574697
R2456 VGND.n431 VGND.n430 0.0574697
R2457 VGND.n606 VGND.n403 0.0574697
R2458 VGND.n490 VGND.n480 0.0574697
R2459 VGND.n1096 VGND.n137 0.0574697
R2460 VGND.n1113 VGND.n1110 0.0574697
R2461 VGND.n1125 VGND.n1124 0.0574697
R2462 VGND.n1158 VGND.n116 0.0574697
R2463 VGND.n64 VGND.n62 0.0574697
R2464 VGND.n974 VGND.n973 0.0574697
R2465 VGND.n932 VGND.n931 0.0574697
R2466 VGND.n228 VGND 0.047375
R2467 VGND.n1291 VGND 0.047375
R2468 VGND.n1255 VGND 0.047375
R2469 VGND VGND.n128 0.047375
R2470 VGND.n110 VGND 0.047375
R2471 VGND.n299 VGND.n233 0.0410405
R2472 VGND.n291 VGND.n289 0.0410405
R2473 VGND.n1339 VGND.n9 0.0410405
R2474 VGND.n11 VGND.n4 0.0410405
R2475 VGND.n1005 VGND.n1004 0.0410405
R2476 VGND.n1007 VGND.n1006 0.0410405
R2477 VGND.n453 VGND.n452 0.0410405
R2478 VGND.n455 VGND.n454 0.0410405
R2479 VGND.n816 VGND.n170 0.0410405
R2480 VGND.n1212 VGND.n1209 0.0410405
R2481 VGND.n1259 VGND.n1210 0.0410405
R2482 VGND.n1300 VGND.n40 0.0410405
R2483 VGND.n1293 VGND.n47 0.0410405
R2484 VGND.n755 VGND.n752 0.0410405
R2485 VGND.n761 VGND.n193 0.0410405
R2486 VGND.n802 VGND.n800 0.0410405
R2487 VGND.n620 VGND.n399 0.0410405
R2488 VGND.n670 VGND.n400 0.0410405
R2489 VGND.n323 VGND.n322 0.0410405
R2490 VGND.n325 VGND.n324 0.0410405
R2491 VGND.n746 VGND.n307 0.0410405
R2492 VGND.n737 VGND.n735 0.0410405
R2493 VGND.n355 VGND.n346 0.0410405
R2494 VGND.n896 VGND.n150 0.0410405
R2495 VGND.n887 VGND.n885 0.0410405
R2496 VGND.n429 VGND.n420 0.0410405
R2497 VGND.n616 VGND.n405 0.0410405
R2498 VGND.n609 VGND.n607 0.0410405
R2499 VGND.n477 VGND.n475 0.0410405
R2500 VGND.n491 VGND.n476 0.0410405
R2501 VGND.n1106 VGND.n139 0.0410405
R2502 VGND.n1099 VGND.n1097 0.0410405
R2503 VGND.n1111 VGND.n132 0.0410405
R2504 VGND.n1126 VGND.n133 0.0410405
R2505 VGND.n853 VGND.n852 0.0410405
R2506 VGND.n1157 VGND.n1156 0.0410405
R2507 VGND.n68 VGND.n61 0.0410405
R2508 VGND.n69 VGND.n65 0.0410405
R2509 VGND.n972 VGND.n922 0.0410405
R2510 VGND.n930 VGND.n924 0.0410405
R2511 VGND.n257 VGND.n31 0.0410405
R2512 VGND.n1308 VGND.n33 0.0410405
R2513 VGND.n333 VGND 0.0382604
R2514 VGND.n762 VGND 0.0369583
R2515 VGND.n1294 VGND 0.0369583
R2516 VGND VGND.n1216 0.0369583
R2517 VGND.n397 VGND 0.0369583
R2518 VGND.n130 VGND 0.0369583
R2519 VGND.n72 VGND 0.0369583
R2520 VGND.n925 VGND 0.0369583
R2521 VGND.n1287 VGND 0.0343542
R2522 VGND VGND.n365 0.0343542
R2523 VGND VGND.n628 0.0343542
R2524 VGND.n543 VGND 0.0343542
R2525 VGND.n1186 VGND 0.0343542
R2526 VGND.n782 VGND 0.0330521
R2527 VGND.n1286 VGND 0.0330521
R2528 VGND.n381 VGND 0.0330521
R2529 VGND.n696 VGND 0.0330521
R2530 VGND VGND.n444 0.0330521
R2531 VGND VGND.n550 0.0330521
R2532 VGND.n871 VGND 0.0330521
R2533 VGND VGND.n50 0.0330521
R2534 VGND VGND.n915 0.0330521
R2535 VGND.n1088 VGND 0.0330521
R2536 VGND VGND.n164 0.0330521
R2537 VGND.n1317 VGND 0.0330521
R2538 VGND.n778 VGND 0.03175
R2539 VGND.n207 VGND 0.03175
R2540 VGND.n1285 VGND 0.03175
R2541 VGND.n1275 VGND 0.03175
R2542 VGND VGND.n551 0.03175
R2543 VGND VGND.n555 0.03175
R2544 VGND.n872 VGND 0.03175
R2545 VGND.n988 VGND 0.03175
R2546 VGND.n1087 VGND 0.03175
R2547 VGND.n1077 VGND 0.03175
R2548 VGND.n1373 VGND 0.03175
R2549 VGND.n35 VGND.n34 0.0292489
R2550 VGND.n891 VGND.n154 0.0292489
R2551 VGND.n886 VGND.n153 0.0292489
R2552 VGND.n900 VGND.n893 0.0292489
R2553 VGND.n902 VGND.n151 0.0292489
R2554 VGND.n351 VGND.n350 0.0292489
R2555 VGND.n353 VGND.n352 0.0292489
R2556 VGND.n806 VGND.n174 0.0292489
R2557 VGND.n801 VGND.n172 0.0292489
R2558 VGND.n812 VGND.n808 0.0292489
R2559 VGND.n814 VGND.n171 0.0292489
R2560 VGND.n430 VGND.n421 0.0292489
R2561 VGND.n423 VGND.n421 0.0292489
R2562 VGND.n1108 VGND.n137 0.0292489
R2563 VGND.n1096 VGND.n136 0.0292489
R2564 VGND.n480 VGND.n479 0.0292489
R2565 VGND.n490 VGND.n489 0.0292489
R2566 VGND.n706 VGND.n705 0.0292489
R2567 VGND.n704 VGND.n703 0.0292489
R2568 VGND.n1302 VGND.n38 0.0292489
R2569 VGND.n46 VGND.n36 0.0292489
R2570 VGND.n1307 VGND.n1306 0.0292489
R2571 VGND.n1125 VGND.n134 0.0292489
R2572 VGND.n1110 VGND.n134 0.0292489
R2573 VGND.n116 VGND.n114 0.0292489
R2574 VGND.n1159 VGND.n1158 0.0292489
R2575 VGND.n1164 VGND.n62 0.0292489
R2576 VGND.n112 VGND.n64 0.0292489
R2577 VGND.n1068 VGND.n1067 0.0292489
R2578 VGND.n1066 VGND.n1065 0.0292489
R2579 VGND.n618 VGND.n403 0.0292489
R2580 VGND.n606 VGND.n402 0.0292489
R2581 VGND.n622 VGND.n401 0.0292489
R2582 VGND.n669 VGND.n668 0.0292489
R2583 VGND.n1215 VGND.n1214 0.0292489
R2584 VGND.n1258 VGND.n1257 0.0292489
R2585 VGND.n1341 VGND.n7 0.0292489
R2586 VGND.n1343 VGND.n5 0.0292489
R2587 VGND.n529 VGND.n528 0.0292489
R2588 VGND.n527 VGND.n526 0.0292489
R2589 VGND.n748 VGND.n305 0.0292489
R2590 VGND.n734 VGND.n303 0.0292489
R2591 VGND.n757 VGND.n750 0.0292489
R2592 VGND.n759 VGND.n229 0.0292489
R2593 VGND.n301 VGND.n231 0.0292489
R2594 VGND.n288 VGND.n230 0.0292489
R2595 VGND.n931 VGND.n923 0.0292489
R2596 VGND.n973 VGND.n923 0.0292489
R2597 VGND VGND.n257 0.027527
R2598 VGND.n1162 VGND 0.0254688
R2599 VGND.n1161 VGND 0.0254688
R2600 VGND.n877 VGND 0.0252396
R2601 VGND.n1134 VGND 0.0252396
R2602 VGND.n754 VGND.n753 0.0239375
R2603 VGND.n1299 VGND.n1298 0.0239375
R2604 VGND.n1262 VGND.n1207 0.0239375
R2605 VGND.n745 VGND.n744 0.0239375
R2606 VGND.n331 VGND.n321 0.0239375
R2607 VGND.n334 VGND.n326 0.0239375
R2608 VGND.n687 VGND 0.0239375
R2609 VGND.n673 VGND.n397 0.0239375
R2610 VGND.n624 VGND.n398 0.0239375
R2611 VGND.n459 VGND.n451 0.0239375
R2612 VGND.n462 VGND.n456 0.0239375
R2613 VGND.n494 VGND.n473 0.0239375
R2614 VGND.n481 VGND.n474 0.0239375
R2615 VGND.n615 VGND.n614 0.0239375
R2616 VGND.n611 VGND.n610 0.0239375
R2617 VGND.n851 VGND.n850 0.0239375
R2618 VGND.n1155 VGND.n118 0.0239375
R2619 VGND.n1129 VGND.n130 0.0239375
R2620 VGND.n1115 VGND.n131 0.0239375
R2621 VGND.n67 VGND.n60 0.0239375
R2622 VGND.n926 VGND.n925 0.0239375
R2623 VGND.n969 VGND.n927 0.0239375
R2624 VGND.n1105 VGND.n1104 0.0239375
R2625 VGND.n1101 VGND.n1100 0.0239375
R2626 VGND.n1014 VGND.n1003 0.0239375
R2627 VGND.n1017 VGND.n1008 0.0239375
R2628 VGND.n298 VGND.n297 0.0239375
R2629 VGND.n293 VGND.n292 0.0239375
R2630 VGND.n1311 VGND.n30 0.0239375
R2631 VGND.n32 VGND.n26 0.0239375
R2632 VGND.n1338 VGND.n1337 0.0239375
R2633 VGND.n10 VGND.n3 0.0239375
R2634 VGND.n795 VGND 0.0226354
R2635 VGND.n783 VGND 0.0226354
R2636 VGND.n781 VGND 0.0226354
R2637 VGND.n763 VGND 0.0226354
R2638 VGND.n221 VGND 0.0226354
R2639 VGND.n218 VGND 0.0226354
R2640 VGND.n1295 VGND 0.0226354
R2641 VGND.n1290 VGND 0.0226354
R2642 VGND.n1281 VGND 0.0226354
R2643 VGND.n1276 VGND 0.0226354
R2644 VGND.n1270 VGND 0.0226354
R2645 VGND VGND.n1208 0.0226354
R2646 VGND.n1254 VGND 0.0226354
R2647 VGND.n1241 VGND 0.0226354
R2648 VGND.n357 VGND 0.0226354
R2649 VGND.n739 VGND 0.0226354
R2650 VGND VGND.n311 0.0226354
R2651 VGND.n713 VGND 0.0226354
R2652 VGND VGND.n331 0.0226354
R2653 VGND VGND.n327 0.0226354
R2654 VGND VGND.n386 0.0226354
R2655 VGND.n681 VGND 0.0226354
R2656 VGND.n661 VGND 0.0226354
R2657 VGND.n653 VGND 0.0226354
R2658 VGND VGND.n631 0.0226354
R2659 VGND VGND.n635 0.0226354
R2660 VGND.n426 VGND 0.0226354
R2661 VGND VGND.n443 0.0226354
R2662 VGND.n539 VGND 0.0226354
R2663 VGND.n515 VGND 0.0226354
R2664 VGND.n511 VGND 0.0226354
R2665 VGND.n486 VGND 0.0226354
R2666 VGND.n482 VGND 0.0226354
R2667 VGND VGND.n565 0.0226354
R2668 VGND.n590 VGND 0.0226354
R2669 VGND.n158 VGND 0.0226354
R2670 VGND.n850 VGND 0.0226354
R2671 VGND.n1137 VGND 0.0226354
R2672 VGND.n1116 VGND 0.0226354
R2673 VGND.n1170 VGND 0.0226354
R2674 VGND.n102 VGND 0.0226354
R2675 VGND.n99 VGND 0.0226354
R2676 VGND.n85 VGND 0.0226354
R2677 VGND.n894 VGND 0.0226354
R2678 VGND VGND.n914 0.0226354
R2679 VGND.n959 VGND 0.0226354
R2680 VGND.n949 VGND 0.0226354
R2681 VGND.n1092 VGND 0.0226354
R2682 VGND VGND.n995 0.0226354
R2683 VGND VGND.n1009 0.0226354
R2684 VGND.n1056 VGND 0.0226354
R2685 VGND.n1048 VGND 0.0226354
R2686 VGND VGND.n1026 0.0226354
R2687 VGND VGND.n1030 0.0226354
R2688 VGND.n818 VGND 0.0226354
R2689 VGND.n832 VGND 0.0226354
R2690 VGND.n247 VGND 0.0226354
R2691 VGND VGND.n251 0.0226354
R2692 VGND.n270 VGND 0.0226354
R2693 VGND.n262 VGND 0.0226354
R2694 VGND.n261 VGND 0.0226354
R2695 VGND VGND.n1320 0.0226354
R2696 VGND VGND.n1325 0.0226354
R2697 VGND.n1333 VGND 0.0226354
R2698 VGND.n1379 VGND 0.0226354
R2699 VGND.n1370 VGND 0.0226354
R2700 VGND.n1355 VGND 0.0226354
R2701 VGND VGND.n202 0.0213333
R2702 VGND.n1240 VGND 0.0213333
R2703 VGND VGND.n572 0.0213333
R2704 VGND VGND.n1021 0.0213333
R2705 VGND.n73 VGND 0.0200312
R2706 VGND.n770 VGND.n187 0.0135208
R2707 VGND.n228 VGND.n227 0.0135208
R2708 VGND.n206 VGND.n39 0.0135208
R2709 VGND.n1291 VGND.n1290 0.0135208
R2710 VGND.n1211 VGND.n1205 0.0135208
R2711 VGND.n1255 VGND.n1254 0.0135208
R2712 VGND.n370 VGND.n306 0.0135208
R2713 VGND.n732 VGND.n731 0.0135208
R2714 VGND.n709 VGND.n708 0.0135208
R2715 VGND.n701 VGND.n700 0.0135208
R2716 VGND.n676 VGND.n394 0.0135208
R2717 VGND.n666 VGND.n665 0.0135208
R2718 VGND.n532 VGND.n531 0.0135208
R2719 VGND.n524 VGND.n523 0.0135208
R2720 VGND.n498 VGND.n471 0.0135208
R2721 VGND.n487 VGND.n486 0.0135208
R2722 VGND.n566 VGND.n404 0.0135208
R2723 VGND.n604 VGND.n603 0.0135208
R2724 VGND.n883 VGND.n882 0.0135208
R2725 VGND.n856 VGND.n855 0.0135208
R2726 VGND.n1154 VGND.n1153 0.0135208
R2727 VGND.n1132 VGND.n128 0.0135208
R2728 VGND.n1122 VGND.n1121 0.0135208
R2729 VGND.n1167 VGND.n1166 0.0135208
R2730 VGND.n110 VGND.n109 0.0135208
R2731 VGND.n977 VGND.n976 0.0135208
R2732 VGND.n966 VGND.n934 0.0135208
R2733 VGND.n943 VGND.n138 0.0135208
R2734 VGND.n1094 VGND.n1093 0.0135208
R2735 VGND.n1071 VGND.n1070 0.0135208
R2736 VGND.n1063 VGND.n1062 0.0135208
R2737 VGND.n823 VGND.n168 0.0135208
R2738 VGND.n235 VGND.n232 0.0135208
R2739 VGND.n286 VGND.n285 0.0135208
R2740 VGND.n260 VGND.n259 0.0135208
R2741 VGND.n1315 VGND.n25 0.0135208
R2742 VGND.n14 VGND.n8 0.0135208
R2743 VGND.n1346 VGND.n1345 0.0135208
R2744 VGND VGND.n394 0.00961458
R2745 VGND.n976 VGND 0.00961458
R2746 VGND.n892 VGND 0.00755
R2747 VGND.n1114 VGND 0.00755
R2748 VGND.n1163 VGND 0.00755
R2749 VGND VGND.n1160 0.00755
R2750 VGND VGND.n72 0.00440625
R2751 VGND.n799 VGND 0.00180208
R2752 VGND VGND.n762 0.00180208
R2753 VGND VGND.n1294 0.00180208
R2754 VGND.n1216 VGND 0.00180208
R2755 VGND VGND.n356 0.00180208
R2756 VGND VGND.n738 0.00180208
R2757 VGND VGND.n419 0.00180208
R2758 VGND.n884 VGND 0.00180208
R2759 VGND VGND.n149 0.00180208
R2760 VGND VGND.n817 0.00180208
R2761 VPWR.n877 VPWR.t49 836.124
R2762 VPWR.n433 VPWR.t311 835.927
R2763 VPWR.n786 VPWR.t43 832.876
R2764 VPWR VPWR.t174 820.76
R2765 VPWR VPWR.t119 820.76
R2766 VPWR.t101 VPWR 820.76
R2767 VPWR.n95 VPWR.t159 812.141
R2768 VPWR.n709 VPWR.t175 812.141
R2769 VPWR.n732 VPWR.t120 812.141
R2770 VPWR.n451 VPWR.t208 812.141
R2771 VPWR.n493 VPWR.t102 812.141
R2772 VPWR.n553 VPWR.t209 812.014
R2773 VPWR.n1008 VPWR.t223 811.918
R2774 VPWR.n689 VPWR.t156 811.918
R2775 VPWR.n676 VPWR.t235 811.918
R2776 VPWR.n760 VPWR.t256 809.183
R2777 VPWR.n358 VPWR.t245 807.481
R2778 VPWR.n922 VPWR.t183 806.484
R2779 VPWR.n813 VPWR.t238 804.731
R2780 VPWR.n349 VPWR.t190 804.731
R2781 VPWR.n352 VPWR.t250 804.731
R2782 VPWR.n39 VPWR.t193 804.731
R2783 VPWR.n367 VPWR.t192 804.731
R2784 VPWR.n366 VPWR.t246 804.731
R2785 VPWR.n345 VPWR.t99 804.731
R2786 VPWR.n1082 VPWR.t229 804.731
R2787 VPWR.n1085 VPWR.t130 804.731
R2788 VPWR.n896 VPWR.t240 804.731
R2789 VPWR.n899 VPWR.t136 804.731
R2790 VPWR.n86 VPWR.t224 804.731
R2791 VPWR.n974 VPWR.t158 804.731
R2792 VPWR.n312 VPWR.t215 804.731
R2793 VPWR.n314 VPWR.t162 804.731
R2794 VPWR.n946 VPWR.t214 804.731
R2795 VPWR.n941 VPWR.t161 804.731
R2796 VPWR.n325 VPWR.t112 804.731
R2797 VPWR.n327 VPWR.t184 804.731
R2798 VPWR.n923 VPWR.t111 804.731
R2799 VPWR.t164 VPWR.n906 804.731
R2800 VPWR.n1035 VPWR.t147 804.731
R2801 VPWR.n1049 VPWR.t124 804.731
R2802 VPWR.n1052 VPWR.t173 804.731
R2803 VPWR.n419 VPWR.t127 804.731
R2804 VPWR.n422 VPWR.t178 804.731
R2805 VPWR.n727 VPWR.t176 804.731
R2806 VPWR.n695 VPWR.t155 804.731
R2807 VPWR.n759 VPWR.t121 804.731
R2808 VPWR.n439 VPWR.t255 804.731
R2809 VPWR.t211 VPWR.n429 804.731
R2810 VPWR.n818 VPWR.t168 804.731
R2811 VPWR.n821 VPWR.t219 804.731
R2812 VPWR.n465 VPWR.t171 804.731
R2813 VPWR.n468 VPWR.t221 804.731
R2814 VPWR.n582 VPWR.t150 804.731
R2815 VPWR.n555 VPWR.t149 804.731
R2816 VPWR.n678 VPWR.t103 804.731
R2817 VPWR.n520 VPWR.t234 804.731
R2818 VPWR.t137 VPWR.n488 804.731
R2819 VPWR.n607 VPWR.t217 804.731
R2820 VPWR.n610 VPWR.t109 804.731
R2821 VPWR.n20 VPWR.t253 804.731
R2822 VPWR.n10 VPWR.t252 804.731
R2823 VPWR.n118 VPWR.t133 804.731
R2824 VPWR.n155 VPWR.t199 804.731
R2825 VPWR.n159 VPWR.t207 804.731
R2826 VPWR.n235 VPWR.t232 804.731
R2827 VPWR.n238 VPWR.t248 804.731
R2828 VPWR.t99 VPWR.n344 751.692
R2829 VPWR.n907 VPWR.t164 751.692
R2830 VPWR.n430 VPWR.t211 751.692
R2831 VPWR.n489 VPWR.t137 751.692
R2832 VPWR.t238 VPWR.n812 725.173
R2833 VPWR.t190 VPWR.n348 725.173
R2834 VPWR.t250 VPWR.n351 725.173
R2835 VPWR.t229 VPWR.n1081 725.173
R2836 VPWR.t130 VPWR.n1084 725.173
R2837 VPWR.t240 VPWR.n895 725.173
R2838 VPWR.t136 VPWR.n898 725.173
R2839 VPWR.t147 VPWR.n1034 725.173
R2840 VPWR.t124 VPWR.n1048 725.173
R2841 VPWR.t173 VPWR.n1051 725.173
R2842 VPWR.t127 VPWR.n418 725.173
R2843 VPWR.t178 VPWR.n421 725.173
R2844 VPWR.t168 VPWR.n817 725.173
R2845 VPWR.t219 VPWR.n820 725.173
R2846 VPWR.t171 VPWR.n464 725.173
R2847 VPWR.t221 VPWR.n467 725.173
R2848 VPWR.t217 VPWR.n606 725.173
R2849 VPWR.t109 VPWR.n609 725.173
R2850 VPWR.t133 VPWR.n117 725.173
R2851 VPWR.t199 VPWR.n154 725.173
R2852 VPWR.t207 VPWR.n158 725.173
R2853 VPWR.t232 VPWR.n234 725.173
R2854 VPWR.t248 VPWR.n237 725.173
R2855 VPWR.t154 VPWR 723.41
R2856 VPWR.t254 VPWR 723.41
R2857 VPWR VPWR.t233 723.41
R2858 VPWR.n1109 VPWR.n61 721.278
R2859 VPWR.n1101 VPWR.n69 721.278
R2860 VPWR.n793 VPWR.n792 721.278
R2861 VPWR.n92 VPWR.n91 713.462
R2862 VPWR.n1115 VPWR.t33 700.506
R2863 VPWR.n1095 VPWR.t367 700.506
R2864 VPWR.n1103 VPWR.t20 698.091
R2865 VPWR.n1116 VPWR.t390 669.491
R2866 VPWR.n62 VPWR.t302 669.491
R2867 VPWR.n840 VPWR.t483 665.307
R2868 VPWR.n1103 VPWR.n65 615.659
R2869 VPWR.n89 VPWR.n88 609.847
R2870 VPWR.n853 VPWR.n791 607.155
R2871 VPWR.n76 VPWR.n75 604.076
R2872 VPWR.n616 VPWR.n602 604.076
R2873 VPWR.n616 VPWR.n603 604.076
R2874 VPWR.n143 VPWR.n110 604.076
R2875 VPWR.n1166 VPWR.n23 604.076
R2876 VPWR.n281 VPWR.n199 604.076
R2877 VPWR.n244 VPWR.n230 604.076
R2878 VPWR.n244 VPWR.n231 604.076
R2879 VPWR.n1026 VPWR.n1025 603.859
R2880 VPWR.n799 VPWR.n798 603.859
R2881 VPWR.n56 VPWR.n55 603.38
R2882 VPWR.n846 VPWR.n795 603.38
R2883 VPWR.n633 VPWR.n584 603.263
R2884 VPWR.n213 VPWR.n212 603.106
R2885 VPWR.n1037 VPWR.n1036 599.808
R2886 VPWR.n8 VPWR.n7 599.808
R2887 VPWR.n15 VPWR.n14 599.808
R2888 VPWR.n168 VPWR.n151 599.808
R2889 VPWR.n204 VPWR.n203 599.808
R2890 VPWR.n268 VPWR.n207 599.808
R2891 VPWR.t185 VPWR 568.994
R2892 VPWR.t151 VPWR.t134 540.46
R2893 VPWR.t200 VPWR.t125 540.46
R2894 VPWR.t113 VPWR 515.284
R2895 VPWR VPWR.t182 511.926
R2896 VPWR VPWR.t160 511.926
R2897 VPWR VPWR.t203 511.926
R2898 VPWR VPWR.t188 493.464
R2899 VPWR.n893 VPWR 491.784
R2900 VPWR.t142 VPWR.t60 466.608
R2901 VPWR.t182 VPWR.t110 463.252
R2902 VPWR.t160 VPWR.t213 463.252
R2903 VPWR.t203 VPWR.t148 463.252
R2904 VPWR.t110 VPWR 414.577
R2905 VPWR.t213 VPWR 414.577
R2906 VPWR.t225 VPWR 414.577
R2907 VPWR VPWR.t113 414.577
R2908 VPWR.t295 VPWR.t107 404.505
R2909 VPWR.t341 VPWR.t197 404.505
R2910 VPWR.t322 VPWR.t230 404.505
R2911 VPWR.n902 VPWR.t153 396.406
R2912 VPWR.n425 VPWR.t202 396.406
R2913 VPWR.n665 VPWR.t144 396.406
R2914 VPWR.t443 VPWR.t128 396.113
R2915 VPWR.n901 VPWR.t152 391.005
R2916 VPWR.n424 VPWR.t201 391.005
R2917 VPWR.n456 VPWR.t143 391.005
R2918 VPWR.n696 VPWR.t212 390.913
R2919 VPWR.n525 VPWR.t138 390.913
R2920 VPWR.n342 VPWR.t100 389.526
R2921 VPWR.n333 VPWR.t165 389.195
R2922 VPWR.n396 VPWR.t186 388.656
R2923 VPWR.n366 VPWR.t187 388.656
R2924 VPWR.n43 VPWR.t180 388.656
R2925 VPWR.n1129 VPWR.t181 388.656
R2926 VPWR.n777 VPWR.t140 388.656
R2927 VPWR.n861 VPWR.t141 388.656
R2928 VPWR.n800 VPWR.t195 388.656
R2929 VPWR.n815 VPWR.t196 388.656
R2930 VPWR.n473 VPWR.t242 388.656
R2931 VPWR.n460 VPWR.t243 388.656
R2932 VPWR.n535 VPWR.t114 388.656
R2933 VPWR.n527 VPWR.t115 388.656
R2934 VPWR.n162 VPWR.t105 388.656
R2935 VPWR.n169 VPWR.t106 388.656
R2936 VPWR.n984 VPWR.t226 388.656
R2937 VPWR.n1003 VPWR.t227 388.656
R2938 VPWR.n644 VPWR.t205 388.656
R2939 VPWR.n654 VPWR.t204 385.026
R2940 VPWR.n50 VPWR.t117 381.443
R2941 VPWR.n1118 VPWR.t118 381.443
R2942 VPWR.n811 VPWR.t237 380.193
R2943 VPWR.n347 VPWR.t189 380.193
R2944 VPWR.n350 VPWR.t249 380.193
R2945 VPWR.n1080 VPWR.t228 380.193
R2946 VPWR.n1083 VPWR.t129 380.193
R2947 VPWR.n894 VPWR.t239 380.193
R2948 VPWR.n897 VPWR.t135 380.193
R2949 VPWR.n1033 VPWR.t146 380.193
R2950 VPWR.n1047 VPWR.t123 380.193
R2951 VPWR.n1050 VPWR.t172 380.193
R2952 VPWR.n417 VPWR.t126 380.193
R2953 VPWR.n420 VPWR.t177 380.193
R2954 VPWR.n816 VPWR.t167 380.193
R2955 VPWR.n819 VPWR.t218 380.193
R2956 VPWR.n463 VPWR.t170 380.193
R2957 VPWR.n466 VPWR.t220 380.193
R2958 VPWR.n605 VPWR.t216 380.193
R2959 VPWR.n608 VPWR.t108 380.193
R2960 VPWR.n116 VPWR.t132 380.193
R2961 VPWR.n153 VPWR.t198 380.193
R2962 VPWR.n157 VPWR.t206 380.193
R2963 VPWR.n233 VPWR.t231 380.193
R2964 VPWR.n236 VPWR.t247 380.193
R2965 VPWR VPWR.t244 360.866
R2966 VPWR.n1088 VPWR.t416 344.06
R2967 VPWR.n604 VPWR.t296 344.06
R2968 VPWR.n256 VPWR.t280 344.06
R2969 VPWR.n232 VPWR.t455 344.06
R2970 VPWR.n604 VPWR.t437 344.06
R2971 VPWR.n109 VPWR.t3 344.06
R2972 VPWR.n6 VPWR.t93 344.06
R2973 VPWR.n232 VPWR.t323 344.06
R2974 VPWR.n1037 VPWR.t408 340.243
R2975 VPWR.n581 VPWR.t276 340.243
R2976 VPWR.n161 VPWR.t342 340.243
R2977 VPWR.n269 VPWR.t264 340.243
R2978 VPWR.n1179 VPWR.t321 340.241
R2979 VPWR.n19 VPWR.t467 340.241
R2980 VPWR.n201 VPWR.t348 340.241
R2981 VPWR.n209 VPWR.t71 340.241
R2982 VPWR.n881 VPWR 339.046
R2983 VPWR.n550 VPWR 339.046
R2984 VPWR.n633 VPWR.t487 337.95
R2985 VPWR VPWR.t169 337.368
R2986 VPWR.n1089 VPWR.n1079 317.103
R2987 VPWR.n1110 VPWR.n59 315.406
R2988 VPWR.n1102 VPWR.n66 315.406
R2989 VPWR.n120 VPWR.n119 313.575
R2990 VPWR.n359 VPWR.t539 313.42
R2991 VPWR.n878 VPWR.n765 312.827
R2992 VPWR.n142 VPWR.n113 312.053
R2993 VPWR.n22 VPWR.n21 312.053
R2994 VPWR.n187 VPWR.n186 312.053
R2995 VPWR.n282 VPWR.n198 312.053
R2996 VPWR.n790 VPWR.n789 312.051
R2997 VPWR.n108 VPWR.n107 312.051
R2998 VPWR.n213 VPWR.n211 312.051
R2999 VPWR.n1094 VPWR.n74 311.659
R3000 VPWR.n1058 VPWR.n1032 311.659
R3001 VPWR.n586 VPWR.n585 311.659
R3002 VPWR.n590 VPWR.n589 311.659
R3003 VPWR.n217 VPWR.n216 311.659
R3004 VPWR.n590 VPWR.n588 311.659
R3005 VPWR.n141 VPWR.n114 311.659
R3006 VPWR.n135 VPWR.n123 311.659
R3007 VPWR.n283 VPWR.n188 311.659
R3008 VPWR.n217 VPWR.n215 311.659
R3009 VPWR.n1123 VPWR.n49 311.519
R3010 VPWR.n45 VPWR.n42 309.519
R3011 VPWR.n379 VPWR.n369 309.517
R3012 VPWR.n36 VPWR.n35 309.517
R3013 VPWR.t244 VPWR.t185 308.834
R3014 VPWR.t157 VPWR.t225 308.834
R3015 VPWR.n639 VPWR.n580 308.755
R3016 VPWR.n671 VPWR.n452 308.755
R3017 VPWR.n475 VPWR.n462 308.755
R3018 VPWR.n94 VPWR.n93 308.755
R3019 VPWR.n149 VPWR.n148 308.151
R3020 VPWR.n276 VPWR.n202 308.151
R3021 VPWR.n262 VPWR.n210 308.151
R3022 VPWR.n1185 VPWR.n11 308.149
R3023 VPWR.n1173 VPWR.n17 308.149
R3024 VPWR.n271 VPWR.n206 308.149
R3025 VPWR.n370 VPWR.t502 306.735
R3026 VPWR.n331 VPWR.t515 306.735
R3027 VPWR.n929 VPWR.t527 306.735
R3028 VPWR.n318 VPWR.t521 306.735
R3029 VPWR.n962 VPWR.t494 306.735
R3030 VPWR.n310 VPWR.t522 306.735
R3031 VPWR.n1014 VPWR.t546 306.735
R3032 VPWR.n747 VPWR.t541 306.735
R3033 VPWR.n437 VPWR.t536 306.735
R3034 VPWR.n715 VPWR.t516 306.735
R3035 VPWR.n693 VPWR.t514 306.735
R3036 VPWR.n577 VPWR.t513 306.735
R3037 VPWR.n495 VPWR.t530 306.735
R3038 VPWR.n514 VPWR.t547 306.735
R3039 VPWR.n455 VPWR.t497 306.735
R3040 VPWR.n12 VPWR.t533 306.735
R3041 VPWR.n774 VPWR.n767 304.731
R3042 VPWR.n859 VPWR.n858 304.731
R3043 VPWR.n774 VPWR.n773 295.255
R3044 VPWR.n859 VPWR.n788 295.255
R3045 VPWR VPWR.t380 290.372
R3046 VPWR VPWR.t478 285.337
R3047 VPWR VPWR.t122 280.3
R3048 VPWR VPWR.t166 280.3
R3049 VPWR.t429 VPWR 271.909
R3050 VPWR VPWR.t98 260.159
R3051 VPWR VPWR.t151 260.159
R3052 VPWR VPWR.t200 260.159
R3053 VPWR VPWR.t142 260.159
R3054 VPWR VPWR.t241 256.803
R3055 VPWR.n812 VPWR.t544 245.667
R3056 VPWR.n348 VPWR.t509 245.667
R3057 VPWR.n351 VPWR.t537 245.667
R3058 VPWR.n1081 VPWR.t498 245.667
R3059 VPWR.n1084 VPWR.t520 245.667
R3060 VPWR.n895 VPWR.t496 245.667
R3061 VPWR.n898 VPWR.t519 245.667
R3062 VPWR.n1034 VPWR.t528 245.667
R3063 VPWR.n1048 VPWR.t535 245.667
R3064 VPWR.n1051 VPWR.t503 245.667
R3065 VPWR.n418 VPWR.t534 245.667
R3066 VPWR.n421 VPWR.t505 245.667
R3067 VPWR.n817 VPWR.t517 245.667
R3068 VPWR.n820 VPWR.t493 245.667
R3069 VPWR.n464 VPWR.t504 245.667
R3070 VPWR.n467 VPWR.t492 245.667
R3071 VPWR.n606 VPWR.t491 245.667
R3072 VPWR.n609 VPWR.t532 245.667
R3073 VPWR.n117 VPWR.t529 245.667
R3074 VPWR.n154 VPWR.t507 245.667
R3075 VPWR.n158 VPWR.t500 245.667
R3076 VPWR.n234 VPWR.t495 245.667
R3077 VPWR.n237 VPWR.t538 245.667
R3078 VPWR.n120 VPWR.t383 245.636
R3079 VPWR.n52 VPWR.t525 242.282
R3080 VPWR.t191 VPWR.t38 241.696
R3081 VPWR.t423 VPWR.t394 236.661
R3082 VPWR.t194 VPWR.t236 231.625
R3083 VPWR VPWR.t275 221.555
R3084 VPWR.t320 VPWR 221.555
R3085 VPWR.t466 VPWR 221.555
R3086 VPWR.n373 VPWR.n372 219.787
R3087 VPWR.n1141 VPWR.n38 219.787
R3088 VPWR.n1130 VPWR.n46 219.787
R3089 VPWR.n344 VPWR.t545 214.906
R3090 VPWR.n880 VPWR.n879 213.119
R3091 VPWR.n909 VPWR.n893 211.137
R3092 VPWR.n44 VPWR.t512 210.964
R3093 VPWR.n901 VPWR.t526 210.964
R3094 VPWR.n424 VPWR.t508 210.964
R3095 VPWR.n474 VPWR.t540 210.964
R3096 VPWR.n456 VPWR.t518 210.964
R3097 VPWR.n152 VPWR.t542 210.964
R3098 VPWR.n1124 VPWR.n48 209.368
R3099 VPWR.n405 VPWR.n341 209.368
R3100 VPWR.n979 VPWR.n311 209.368
R3101 VPWR.n882 VPWR.n881 209.368
R3102 VPWR.n660 VPWR.n550 209.368
R3103 VPWR.n179 VPWR.n178 209.368
R3104 VPWR VPWR.t157 206.45
R3105 VPWR VPWR.t56 206.45
R3106 VPWR VPWR.t11 206.45
R3107 VPWR VPWR.t257 206.45
R3108 VPWR.t430 VPWR 196.379
R3109 VPWR.t128 VPWR 182.952
R3110 VPWR.t122 VPWR 182.952
R3111 VPWR.t236 VPWR 182.952
R3112 VPWR.t166 VPWR 182.952
R3113 VPWR.t107 VPWR 182.952
R3114 VPWR.t230 VPWR 182.952
R3115 VPWR.n341 VPWR 179.595
R3116 VPWR.t380 VPWR.t299 179.595
R3117 VPWR.t38 VPWR.t387 179.595
R3118 VPWR.t52 VPWR.t440 179.595
R3119 VPWR.n311 VPWR 179.595
R3120 VPWR VPWR.n549 179.595
R3121 VPWR.n180 VPWR 179.595
R3122 VPWR.t470 VPWR.t385 162.81
R3123 VPWR.t484 VPWR.t54 162.81
R3124 VPWR.t478 VPWR.t307 162.81
R3125 VPWR.t80 VPWR.t480 162.81
R3126 VPWR.t391 VPWR 161.131
R3127 VPWR.t376 VPWR.t297 161.131
R3128 VPWR.t359 VPWR.t90 161.131
R3129 VPWR.t58 VPWR.t318 161.131
R3130 VPWR.t332 VPWR.t488 161.131
R3131 VPWR.t445 VPWR.t265 161.131
R3132 VPWR.t433 VPWR.t281 161.131
R3133 VPWR.t287 VPWR.t324 161.131
R3134 VPWR.t372 VPWR.t23 159.452
R3135 VPWR.t50 VPWR.t14 159.452
R3136 VPWR.t139 VPWR.t42 157.774
R3137 VPWR.t396 VPWR.t447 156.095
R3138 VPWR.t174 VPWR.t154 154.417
R3139 VPWR.t119 VPWR.t254 154.417
R3140 VPWR.t233 VPWR.t101 154.417
R3141 VPWR.t385 VPWR 152.739
R3142 VPWR.t54 VPWR 152.739
R3143 VPWR.t474 VPWR 152.739
R3144 VPWR.t78 VPWR.t427 152.739
R3145 VPWR.t458 VPWR.t72 152.739
R3146 VPWR.t11 VPWR.t222 151.06
R3147 VPWR.t301 VPWR.t19 147.703
R3148 VPWR.t56 VPWR.t62 147.703
R3149 VPWR.t449 VPWR.t46 147.703
R3150 VPWR.t411 VPWR.t40 147.703
R3151 VPWR.t60 VPWR.t303 147.703
R3152 VPWR.t257 VPWR.t74 147.703
R3153 VPWR.t8 VPWR.t431 147.703
R3154 VPWR.t413 VPWR.t415 144.346
R3155 VPWR.t403 VPWR.t405 144.346
R3156 VPWR.t269 VPWR.t271 144.346
R3157 VPWR.t297 VPWR.t291 144.346
R3158 VPWR.t291 VPWR.t293 144.346
R3159 VPWR.t293 VPWR.t295 144.346
R3160 VPWR.t339 VPWR.t337 144.346
R3161 VPWR.t88 VPWR.t86 144.346
R3162 VPWR.t90 VPWR.t88 144.346
R3163 VPWR.t316 VPWR.t314 144.346
R3164 VPWR.t318 VPWR.t316 144.346
R3165 VPWR.t2 VPWR.t6 144.346
R3166 VPWR.t343 VPWR.t349 144.346
R3167 VPWR.t64 VPWR.t66 144.346
R3168 VPWR.t324 VPWR.t326 144.346
R3169 VPWR.t326 VPWR.t328 144.346
R3170 VPWR.t328 VPWR.t322 144.346
R3171 VPWR.t84 VPWR.t285 142.668
R3172 VPWR.t299 VPWR.t470 140.989
R3173 VPWR.t387 VPWR.t484 140.989
R3174 VPWR.t289 VPWR.t363 140.989
R3175 VPWR.t267 VPWR.t21 140.989
R3176 VPWR.t447 VPWR.t472 140.989
R3177 VPWR.t42 VPWR.t44 140.989
R3178 VPWR.t334 VPWR.t430 140.989
R3179 VPWR.t351 VPWR.t261 140.989
R3180 VPWR VPWR.t52 139.311
R3181 VPWR.t442 VPWR.t76 139.311
R3182 VPWR.t464 VPWR.t277 139.311
R3183 VPWR.t305 VPWR.t0 139.311
R3184 VPWR.t345 VPWR.t399 139.311
R3185 VPWR.t355 VPWR.t279 139.311
R3186 VPWR.t451 VPWR.t30 137.633
R3187 VPWR.t425 VPWR.t34 137.633
R3188 VPWR.t104 VPWR.t341 135.954
R3189 VPWR.t251 VPWR.t320 135.954
R3190 VPWR.t26 VPWR.t96 132.597
R3191 VPWR.t28 VPWR.t421 132.597
R3192 VPWR.t419 VPWR.t24 132.597
R3193 VPWR.n810 VPWR.t511 129.344
R3194 VPWR.n985 VPWR.t543 129.344
R3195 VPWR.n867 VPWR.t531 129.344
R3196 VPWR.n534 VPWR.t524 129.344
R3197 VPWR VPWR.t334 127.562
R3198 VPWR.t188 VPWR 125.883
R3199 VPWR.n341 VPWR 125.883
R3200 VPWR.t134 VPWR 125.883
R3201 VPWR VPWR.n311 125.883
R3202 VPWR VPWR.t393 125.883
R3203 VPWR.t125 VPWR 125.883
R3204 VPWR.t169 VPWR 125.883
R3205 VPWR.n549 VPWR 125.883
R3206 VPWR.n550 VPWR 125.883
R3207 VPWR.t197 VPWR 125.883
R3208 VPWR VPWR.t2 125.883
R3209 VPWR.t407 VPWR 124.206
R3210 VPWR.n180 VPWR 124.206
R3211 VPWR.t68 VPWR.t263 124.206
R3212 VPWR.t362 VPWR.t439 120.849
R3213 VPWR.t16 VPWR.t429 120.849
R3214 VPWR.t279 VPWR 120.849
R3215 VPWR.t486 VPWR.t273 119.171
R3216 VPWR.n907 VPWR.t506 118.853
R3217 VPWR.n430 VPWR.t499 118.853
R3218 VPWR.t439 VPWR 117.492
R3219 VPWR.n394 VPWR.t510 117.294
R3220 VPWR.t490 VPWR 115.814
R3221 VPWR.t417 VPWR.t365 115.814
R3222 VPWR.t44 VPWR 115.814
R3223 VPWR.t349 VPWR 114.135
R3224 VPWR.t66 VPWR 114.135
R3225 VPWR.t312 VPWR 112.457
R3226 VPWR.n490 VPWR.t523 111.576
R3227 VPWR.n652 VPWR.t501 111.537
R3228 VPWR.t36 VPWR 110.778
R3229 VPWR.t14 VPWR 110.778
R3230 VPWR.t368 VPWR 110.778
R3231 VPWR VPWR.t374 110.778
R3232 VPWR VPWR.t359 110.778
R3233 VPWR VPWR.t58 110.778
R3234 VPWR VPWR.t78 110.778
R3235 VPWR.t19 VPWR 109.1
R3236 VPWR.t366 VPWR 109.1
R3237 VPWR.t62 VPWR 109.1
R3238 VPWR.t472 VPWR 109.1
R3239 VPWR.t74 VPWR 109.1
R3240 VPWR.t431 VPWR 109.1
R3241 VPWR.t384 VPWR 107.421
R3242 VPWR VPWR.t339 107.421
R3243 VPWR VPWR.t382 107.421
R3244 VPWR.n549 VPWR.n548 106.561
R3245 VPWR.n181 VPWR.n180 106.561
R3246 VPWR.t148 VPWR 105.743
R3247 VPWR.t309 VPWR.t370 104.064
R3248 VPWR VPWR.t4 104.064
R3249 VPWR.t389 VPWR 102.385
R3250 VPWR.t10 VPWR.t409 102.385
R3251 VPWR.t378 VPWR 102.385
R3252 VPWR.t401 VPWR 100.707
R3253 VPWR.t179 VPWR.t391 99.0288
R3254 VPWR.t353 VPWR 99.0288
R3255 VPWR.t48 VPWR 99.0288
R3256 VPWR.n1079 VPWR.t25 98.5005
R3257 VPWR VPWR.t468 97.3503
R3258 VPWR.n49 VPWR.t373 96.1553
R3259 VPWR.n59 VPWR.t27 96.1553
R3260 VPWR.n66 VPWR.t29 96.1553
R3261 VPWR.n1025 VPWR.t479 96.1553
R3262 VPWR.n791 VPWR.t81 96.1553
R3263 VPWR.n798 VPWR.t395 96.1553
R3264 VPWR.n48 VPWR.t372 95.6719
R3265 VPWR.n372 VPWR.t386 95.3969
R3266 VPWR.n38 VPWR.t55 95.3969
R3267 VPWR.n46 VPWR.t475 95.3969
R3268 VPWR.t409 VPWR 93.9934
R3269 VPWR.t482 VPWR.t476 93.9934
R3270 VPWR.t265 VPWR 93.9934
R3271 VPWR.t281 VPWR 93.9934
R3272 VPWR.n61 VPWR.t31 93.81
R3273 VPWR.n69 VPWR.t35 93.81
R3274 VPWR.n91 VPWR.t397 93.81
R3275 VPWR.n792 VPWR.t18 93.81
R3276 VPWR.t370 VPWR 92.315
R3277 VPWR.n179 VPWR.t335 88.9581
R3278 VPWR.t275 VPWR 87.2797
R3279 VPWR VPWR.t466 87.2797
R3280 VPWR.t405 VPWR.t145 85.6012
R3281 VPWR.t46 VPWR.t80 85.6012
R3282 VPWR.t398 VPWR.t17 85.6012
R3283 VPWR VPWR.t92 83.9228
R3284 VPWR.n893 VPWR.t163 77.209
R3285 VPWR.n881 VPWR.t210 77.209
R3286 VPWR.t310 VPWR.n880 73.8521
R3287 VPWR.t460 VPWR.t398 73.8521
R3288 VPWR.t382 VPWR.t131 73.8521
R3289 VPWR.t374 VPWR.n179 72.1736
R3290 VPWR.t330 VPWR.n48 68.8168
R3291 VPWR.t394 VPWR.t482 68.8168
R3292 VPWR.t116 VPWR.t490 67.1383
R3293 VPWR.n880 VPWR.t312 67.1383
R3294 VPWR.t480 VPWR.t460 67.1383
R3295 VPWR.t92 VPWR 67.1383
R3296 VPWR.t131 VPWR.t332 67.1383
R3297 VPWR.n55 VPWR.t290 63.3219
R3298 VPWR.n55 VPWR.t364 63.3219
R3299 VPWR.n65 VPWR.t268 63.3219
R3300 VPWR.n65 VPWR.t22 63.3219
R3301 VPWR.n88 VPWR.t448 63.3219
R3302 VPWR.n88 VPWR.t473 63.3219
R3303 VPWR.n795 VPWR.t371 63.3219
R3304 VPWR.n795 VPWR.t424 63.3219
R3305 VPWR.t86 VPWR 60.4245
R3306 VPWR.t82 VPWR.t10 58.7461
R3307 VPWR.t145 VPWR.t407 58.7461
R3308 VPWR VPWR.t330 57.0676
R3309 VPWR VPWR.t13 57.0676
R3310 VPWR VPWR.t269 57.0676
R3311 VPWR.t468 VPWR 57.0676
R3312 VPWR.n653 VPWR.n652 55.5913
R3313 VPWR.t17 VPWR.t309 55.3892
R3314 VPWR.t23 VPWR.t116 53.7107
R3315 VPWR VPWR.t353 53.7107
R3316 VPWR VPWR.t82 53.7107
R3317 VPWR VPWR.t376 53.7107
R3318 VPWR.t72 VPWR 53.7107
R3319 VPWR VPWR.t401 53.7107
R3320 VPWR VPWR.t287 53.7107
R3321 VPWR VPWR.t289 52.0323
R3322 VPWR VPWR.t310 52.0323
R3323 VPWR VPWR.t48 52.0323
R3324 VPWR VPWR.t139 52.0323
R3325 VPWR VPWR.t449 52.0323
R3326 VPWR.t40 VPWR 52.0323
R3327 VPWR.t303 VPWR 52.0323
R3328 VPWR.t488 VPWR 52.0323
R3329 VPWR VPWR.t378 52.0323
R3330 VPWR VPWR.t94 52.0323
R3331 VPWR VPWR.t301 50.3539
R3332 VPWR VPWR.t403 50.3539
R3333 VPWR VPWR.t259 50.3539
R3334 VPWR VPWR.t283 50.3539
R3335 VPWR VPWR.t191 48.6754
R3336 VPWR VPWR.t267 48.6754
R3337 VPWR.t163 VPWR 48.6754
R3338 VPWR.t210 VPWR 48.6754
R3339 VPWR VPWR.t423 48.6754
R3340 VPWR VPWR.t194 48.6754
R3341 VPWR.t98 VPWR 46.997
R3342 VPWR VPWR.t36 46.997
R3343 VPWR.t462 VPWR 46.997
R3344 VPWR VPWR.t357 45.3185
R3345 VPWR VPWR.t32 43.6401
R3346 VPWR VPWR.t366 43.6401
R3347 VPWR VPWR.t368 43.6401
R3348 VPWR.t440 VPWR.t179 41.9616
R3349 VPWR VPWR.t50 41.9616
R3350 VPWR.t6 VPWR 40.2832
R3351 VPWR.n369 VPWR.t300 38.4155
R3352 VPWR.n35 VPWR.t388 38.4155
R3353 VPWR.n42 VPWR.t441 38.4155
R3354 VPWR.n119 VPWR.t489 38.4155
R3355 VPWR.n369 VPWR.t381 37.4305
R3356 VPWR.n35 VPWR.t39 37.4305
R3357 VPWR.n42 VPWR.t53 37.4305
R3358 VPWR.n74 VPWR.t418 37.4305
R3359 VPWR.n1032 VPWR.t410 37.4305
R3360 VPWR.n585 VPWR.t274 37.4305
R3361 VPWR.n588 VPWR.t438 37.4305
R3362 VPWR.n589 VPWR.t298 37.4305
R3363 VPWR.n114 VPWR.t1 37.4305
R3364 VPWR.n123 VPWR.t465 37.4305
R3365 VPWR.n11 VPWR.t91 37.4305
R3366 VPWR.n17 VPWR.t319 37.4305
R3367 VPWR.n148 VPWR.t336 37.4305
R3368 VPWR.n188 VPWR.t346 37.4305
R3369 VPWR.n202 VPWR.t266 37.4305
R3370 VPWR.n206 VPWR.t69 37.4305
R3371 VPWR.n210 VPWR.t282 37.4305
R3372 VPWR.n215 VPWR.t325 37.4305
R3373 VPWR.n216 VPWR.t456 37.4305
R3374 VPWR.t335 VPWR 36.9263
R3375 VPWR.n788 VPWR.t45 36.4455
R3376 VPWR.n765 VPWR.t313 36.4455
R3377 VPWR.n773 VPWR.t51 36.4455
R3378 VPWR.n93 VPWR.t57 36.1587
R3379 VPWR.n93 VPWR.t63 36.1587
R3380 VPWR.n789 VPWR.t450 36.1587
R3381 VPWR.n789 VPWR.t47 36.1587
R3382 VPWR.n580 VPWR.t258 36.1587
R3383 VPWR.n580 VPWR.t75 36.1587
R3384 VPWR.n452 VPWR.t304 36.1587
R3385 VPWR.n452 VPWR.t61 36.1587
R3386 VPWR.n462 VPWR.t41 36.1587
R3387 VPWR.n462 VPWR.t412 36.1587
R3388 VPWR.n113 VPWR.t459 36.1587
R3389 VPWR.n113 VPWR.t306 36.1587
R3390 VPWR.n21 VPWR.t278 36.1587
R3391 VPWR.n21 VPWR.t428 36.1587
R3392 VPWR.n107 VPWR.t379 36.1587
R3393 VPWR.n107 VPWR.t358 36.1587
R3394 VPWR.n186 VPWR.t9 36.1587
R3395 VPWR.n186 VPWR.t432 36.1587
R3396 VPWR.n198 VPWR.t95 36.1587
R3397 VPWR.n198 VPWR.t400 36.1587
R3398 VPWR.n211 VPWR.t85 36.1587
R3399 VPWR.n211 VPWR.t356 36.1587
R3400 VPWR.n1124 VPWR.n47 34.6358
R3401 VPWR.n1100 VPWR.n70 34.6358
R3402 VPWR.n1096 VPWR.n70 34.6358
R3403 VPWR.n628 VPWR.n627 34.6358
R3404 VPWR.n267 VPWR.n208 34.6358
R3405 VPWR.n275 VPWR.n204 34.2593
R3406 VPWR.n848 VPWR.n847 34.0725
R3407 VPWR.n276 VPWR.n275 32.377
R3408 VPWR.n271 VPWR.n270 32.377
R3409 VPWR.n262 VPWR.n261 32.377
R3410 VPWR.n280 VPWR.n201 30.8711
R3411 VPWR.n270 VPWR.n269 30.8711
R3412 VPWR.n209 VPWR.n208 30.8711
R3413 VPWR VPWR.t347 30.2125
R3414 VPWR VPWR.t70 30.2125
R3415 VPWR.t365 VPWR.t419 28.5341
R3416 VPWR.t393 VPWR 28.5341
R3417 VPWR.n61 VPWR.t97 28.5169
R3418 VPWR.n69 VPWR.t422 28.5169
R3419 VPWR.n792 VPWR.t461 28.5169
R3420 VPWR.n178 VPWR.n6 27.8593
R3421 VPWR.n256 VPWR.n255 27.8593
R3422 VPWR.n74 VPWR.t354 27.5805
R3423 VPWR.n75 VPWR.t420 27.5805
R3424 VPWR.n75 VPWR.t414 27.5805
R3425 VPWR.n1032 VPWR.t83 27.5805
R3426 VPWR.n1036 VPWR.t404 27.5805
R3427 VPWR.n1036 VPWR.t406 27.5805
R3428 VPWR.n788 VPWR.t369 27.5805
R3429 VPWR.n765 VPWR.t37 27.5805
R3430 VPWR.n773 VPWR.t15 27.5805
R3431 VPWR.n584 VPWR.t270 27.5805
R3432 VPWR.n584 VPWR.t272 27.5805
R3433 VPWR.n585 VPWR.t77 27.5805
R3434 VPWR.n588 VPWR.t377 27.5805
R3435 VPWR.n589 VPWR.t457 27.5805
R3436 VPWR.n602 VPWR.t435 27.5805
R3437 VPWR.n602 VPWR.t436 27.5805
R3438 VPWR.n603 VPWR.t292 27.5805
R3439 VPWR.n603 VPWR.t294 27.5805
R3440 VPWR.n110 VPWR.t5 27.5805
R3441 VPWR.n110 VPWR.t7 27.5805
R3442 VPWR.n114 VPWR.t73 27.5805
R3443 VPWR.n123 VPWR.t79 27.5805
R3444 VPWR.n23 VPWR.t469 27.5805
R3445 VPWR.n23 VPWR.t463 27.5805
R3446 VPWR.n7 VPWR.t87 27.5805
R3447 VPWR.n7 VPWR.t89 27.5805
R3448 VPWR.n11 VPWR.t360 27.5805
R3449 VPWR.n14 VPWR.t315 27.5805
R3450 VPWR.n14 VPWR.t317 27.5805
R3451 VPWR.n17 VPWR.t59 27.5805
R3452 VPWR.n151 VPWR.t338 27.5805
R3453 VPWR.n151 VPWR.t340 27.5805
R3454 VPWR.n148 VPWR.t375 27.5805
R3455 VPWR.n188 VPWR.t402 27.5805
R3456 VPWR.n199 VPWR.t344 27.5805
R3457 VPWR.n199 VPWR.t350 27.5805
R3458 VPWR.n202 VPWR.t446 27.5805
R3459 VPWR.n206 VPWR.t352 27.5805
R3460 VPWR.n203 VPWR.t260 27.5805
R3461 VPWR.n203 VPWR.t262 27.5805
R3462 VPWR.n207 VPWR.t65 27.5805
R3463 VPWR.n207 VPWR.t67 27.5805
R3464 VPWR.n210 VPWR.t434 27.5805
R3465 VPWR.n212 VPWR.t284 27.5805
R3466 VPWR.n212 VPWR.t286 27.5805
R3467 VPWR.n215 VPWR.t288 27.5805
R3468 VPWR.n216 VPWR.t361 27.5805
R3469 VPWR.n230 VPWR.t327 27.5805
R3470 VPWR.n230 VPWR.t329 27.5805
R3471 VPWR.n231 VPWR.t453 27.5805
R3472 VPWR.n231 VPWR.t454 27.5805
R3473 VPWR.n848 VPWR.n793 27.4829
R3474 VPWR.n1025 VPWR.t308 27.3647
R3475 VPWR.n791 VPWR.t481 27.3647
R3476 VPWR.n798 VPWR.t477 27.3647
R3477 VPWR.n1190 VPWR.n1189 27.0566
R3478 VPWR.n91 VPWR.t12 26.9729
R3479 VPWR.t30 VPWR.t26 26.8556
R3480 VPWR.t96 VPWR.t362 26.8556
R3481 VPWR.t34 VPWR.t28 26.8556
R3482 VPWR.t421 VPWR.t16 26.8556
R3483 VPWR.n1137 VPWR.n1136 26.7859
R3484 VPWR.n1059 VPWR.n1030 26.7859
R3485 VPWR.n49 VPWR.t331 26.5955
R3486 VPWR.n59 VPWR.t452 26.5955
R3487 VPWR.n66 VPWR.t426 26.5955
R3488 VPWR.n119 VPWR.t333 26.5955
R3489 VPWR.n845 VPWR.n796 26.4678
R3490 VPWR.n372 VPWR.t471 26.3637
R3491 VPWR.n38 VPWR.t485 26.3637
R3492 VPWR.n46 VPWR.t392 26.3637
R3493 VPWR.n655 VPWR.n654 26.3341
R3494 VPWR.n1104 VPWR.n62 25.977
R3495 VPWR.n1096 VPWR.n1095 25.977
R3496 VPWR.n1079 VPWR.t444 25.6105
R3497 VPWR.n1109 VPWR.n1108 25.6005
R3498 VPWR.n1101 VPWR.n1100 25.6005
R3499 VPWR.n852 VPWR.n793 25.6005
R3500 VPWR.n616 VPWR.n615 25.6005
R3501 VPWR.n144 VPWR.n143 25.6005
R3502 VPWR.n281 VPWR.n280 25.6005
R3503 VPWR.n244 VPWR.n243 25.6005
R3504 VPWR.n1059 VPWR.n1058 25.224
R3505 VPWR.n628 VPWR.n586 25.224
R3506 VPWR.n627 VPWR.n590 25.224
R3507 VPWR.n141 VPWR.n140 25.224
R3508 VPWR.n136 VPWR.n135 25.224
R3509 VPWR.n284 VPWR.n283 25.224
R3510 VPWR.n255 VPWR.n217 25.224
R3511 VPWR.n1136 VPWR.n40 25.1912
R3512 VPWR.n1128 VPWR.n47 25.1912
R3513 VPWR.t271 VPWR.t486 25.1772
R3514 VPWR.n1111 VPWR.n1110 25.0372
R3515 VPWR.n1103 VPWR.n1102 24.8476
R3516 VPWR.n490 VPWR.n489 24.7622
R3517 VPWR.n1093 VPWR.n76 24.4711
R3518 VPWR.n617 VPWR.n616 24.4711
R3519 VPWR.n245 VPWR.n244 24.4711
R3520 VPWR.n840 VPWR.n839 24.0618
R3521 VPWR.n1108 VPWR.n62 23.7181
R3522 VPWR.n1104 VPWR.n1103 23.7181
R3523 VPWR.n1057 VPWR.n1038 23.7181
R3524 VPWR.n140 VPWR.n121 23.7181
R3525 VPWR.n136 VPWR.n121 23.7181
R3526 VPWR.n182 VPWR.n181 23.7181
R3527 VPWR.n1123 VPWR.n1122 23.6853
R3528 VPWR.t347 VPWR.t445 23.4987
R3529 VPWR.t70 VPWR.t433 23.4987
R3530 VPWR.n170 VPWR.n149 22.9323
R3531 VPWR.n876 VPWR.n767 22.2123
R3532 VPWR.n858 VPWR.n857 22.2123
R3533 VPWR.n857 VPWR.n790 22.2123
R3534 VPWR.n854 VPWR.n790 22.2123
R3535 VPWR.n182 VPWR.n108 22.2123
R3536 VPWR.n284 VPWR.n187 22.2123
R3537 VPWR.n261 VPWR.n213 22.2123
R3538 VPWR.n257 VPWR.n213 22.2123
R3539 VPWR.n799 VPWR.n796 21.8358
R3540 VPWR.t363 VPWR.t451 21.8203
R3541 VPWR.t21 VPWR.t425 21.8203
R3542 VPWR.t273 VPWR.t442 21.8203
R3543 VPWR.n633 VPWR.n632 21.4593
R3544 VPWR.n708 VPWR.n696 20.8436
R3545 VPWR.n525 VPWR.n524 20.8436
R3546 VPWR.n1094 VPWR.n1093 20.7064
R3547 VPWR.n1058 VPWR.n1057 20.7064
R3548 VPWR.n632 VPWR.n586 20.7064
R3549 VPWR.n617 VPWR.n590 20.7064
R3550 VPWR.n245 VPWR.n217 20.7064
R3551 VPWR.t261 VPWR.t68 20.1418
R3552 VPWR.t263 VPWR.t64 20.1418
R3553 VPWR.n653 VPWR.n554 20.0749
R3554 VPWR.n877 VPWR.n876 19.9534
R3555 VPWR.n615 VPWR.n604 19.9534
R3556 VPWR.n144 VPWR.n109 19.9534
R3557 VPWR.n1190 VPWR.n6 19.9534
R3558 VPWR.n257 VPWR.n256 19.9534
R3559 VPWR.n243 VPWR.n232 19.9534
R3560 VPWR.n1167 VPWR.n1166 17.7506
R3561 VPWR.n1116 VPWR.n1115 17.3181
R3562 VPWR.n384 VPWR.n383 17.2339
R3563 VPWR.n1088 VPWR.n1087 16.9417
R3564 VPWR.n611 VPWR.n604 16.9417
R3565 VPWR.n181 VPWR.n109 16.9417
R3566 VPWR.n239 VPWR.n232 16.9417
R3567 VPWR.n634 VPWR.n633 16.2447
R3568 VPWR.n1115 VPWR.n1114 15.5501
R3569 VPWR.n1110 VPWR.n1109 15.4358
R3570 VPWR.n1102 VPWR.n1101 15.4358
R3571 VPWR.n776 VPWR.n774 15.3731
R3572 VPWR.n860 VPWR.n859 15.3731
R3573 VPWR.t307 VPWR 15.1065
R3574 VPWR.n1095 VPWR.n1094 14.3064
R3575 VPWR.n1117 VPWR.n1116 14.2735
R3576 VPWR.n824 VPWR.n823 14.2735
R3577 VPWR.n548 VPWR.n547 14.2735
R3578 VPWR.n472 VPWR.n469 14.2735
R3579 VPWR.n163 VPWR.n160 14.2735
R3580 VPWR.t476 VPWR 13.4281
R3581 VPWR.n1089 VPWR.n76 13.177
R3582 VPWR.n353 VPWR.n346 12.8005
R3583 VPWR.n905 VPWR.n900 12.8005
R3584 VPWR.n1053 VPWR.n1038 12.8005
R3585 VPWR.n428 VPWR.n423 12.8005
R3586 VPWR.n841 VPWR.n799 12.8005
R3587 VPWR.n548 VPWR.n458 12.8005
R3588 VPWR.n143 VPWR.n142 12.0476
R3589 VPWR.n1166 VPWR.n22 12.0476
R3590 VPWR.n282 VPWR.n281 12.0476
R3591 VPWR.t24 VPWR.t413 11.7496
R3592 VPWR.n878 VPWR.n877 11.6711
R3593 VPWR.n909 VPWR.n908 11.3436
R3594 VPWR.n1089 VPWR.n1088 11.2946
R3595 VPWR.n879 VPWR.n878 11.2946
R3596 VPWR.n488 VPWR.n458 10.5744
R3597 VPWR.n1008 VPWR.n1007 9.8812
R3598 VPWR.n731 VPWR.n689 9.8812
R3599 VPWR.n676 VPWR.n675 9.8812
R3600 VPWR.n187 VPWR.n108 9.78874
R3601 VPWR.n405 VPWR.n404 9.73273
R3602 VPWR.n378 VPWR.n377 9.73273
R3603 VPWR.n374 VPWR.n34 9.73273
R3604 VPWR.n1154 VPWR.n34 9.73273
R3605 VPWR.n1154 VPWR.n1153 9.73273
R3606 VPWR.n1143 VPWR.n1142 9.73273
R3607 VPWR.n1009 VPWR.n94 9.73273
R3608 VPWR.n1013 VPWR.n94 9.73273
R3609 VPWR.n1019 VPWR.n1018 9.73273
R3610 VPWR.n1020 VPWR.n1019 9.73273
R3611 VPWR.n1024 VPWR.n1023 9.73273
R3612 VPWR.n1027 VPWR.n1024 9.73273
R3613 VPWR.n672 VPWR.n671 9.73273
R3614 VPWR.n671 VPWR.n453 9.73273
R3615 VPWR.n667 VPWR.n666 9.73273
R3616 VPWR.n664 VPWR.n457 9.73273
R3617 VPWR.n660 VPWR.n457 9.73273
R3618 VPWR.n660 VPWR.n659 9.73273
R3619 VPWR.n659 VPWR.n551 9.73273
R3620 VPWR.n639 VPWR.n578 9.73273
R3621 VPWR.n639 VPWR.n638 9.73273
R3622 VPWR.n1184 VPWR.n1183 9.73273
R3623 VPWR.n1178 VPWR.n1177 9.73273
R3624 VPWR.n1172 VPWR.n1171 9.73273
R3625 VPWR.n1171 VPWR.n18 9.73273
R3626 VPWR.n1007 VPWR.n95 9.65664
R3627 VPWR.n732 VPWR.n731 9.65664
R3628 VPWR.n709 VPWR.n708 9.65664
R3629 VPWR.n524 VPWR.n493 9.65664
R3630 VPWR.n675 VPWR.n451 9.65664
R3631 VPWR.n489 VPWR.n487 9.6005
R3632 VPWR.n1174 VPWR.n15 9.52116
R3633 VPWR.n655 VPWR.n553 9.49016
R3634 VPWR.n854 VPWR.n853 9.41227
R3635 VPWR.n406 VPWR.n405 9.3005
R3636 VPWR.n404 VPWR.n403 9.3005
R3637 VPWR.n398 VPWR.n397 9.3005
R3638 VPWR.n395 VPWR.n363 9.3005
R3639 VPWR.n393 VPWR.n392 9.3005
R3640 VPWR.n391 VPWR.n364 9.3005
R3641 VPWR.n390 VPWR.n389 9.3005
R3642 VPWR.n388 VPWR.n365 9.3005
R3643 VPWR.n387 VPWR.n386 9.3005
R3644 VPWR.n385 VPWR.n384 9.3005
R3645 VPWR.n383 VPWR.n382 9.3005
R3646 VPWR.n381 VPWR.n380 9.3005
R3647 VPWR.n378 VPWR.n368 9.3005
R3648 VPWR.n377 VPWR.n376 9.3005
R3649 VPWR.n375 VPWR.n374 9.3005
R3650 VPWR.n371 VPWR.n34 9.3005
R3651 VPWR.n1155 VPWR.n1154 9.3005
R3652 VPWR.n1153 VPWR.n1152 9.3005
R3653 VPWR.n1144 VPWR.n1143 9.3005
R3654 VPWR.n1142 VPWR.n37 9.3005
R3655 VPWR.n1140 VPWR.n1139 9.3005
R3656 VPWR.n1138 VPWR.n1137 9.3005
R3657 VPWR.n1136 VPWR.n1135 9.3005
R3658 VPWR.n1134 VPWR.n40 9.3005
R3659 VPWR.n1133 VPWR.n1132 9.3005
R3660 VPWR.n1131 VPWR.n41 9.3005
R3661 VPWR.n1128 VPWR.n1127 9.3005
R3662 VPWR.n1126 VPWR.n47 9.3005
R3663 VPWR.n1125 VPWR.n1124 9.3005
R3664 VPWR.n1122 VPWR.n1121 9.3005
R3665 VPWR.n1120 VPWR.n1119 9.3005
R3666 VPWR.n1117 VPWR.n51 9.3005
R3667 VPWR.n1116 VPWR.n53 9.3005
R3668 VPWR.n1115 VPWR.n54 9.3005
R3669 VPWR.n1114 VPWR.n1113 9.3005
R3670 VPWR.n1112 VPWR.n1111 9.3005
R3671 VPWR.n1110 VPWR.n58 9.3005
R3672 VPWR.n1109 VPWR.n60 9.3005
R3673 VPWR.n1108 VPWR.n1107 9.3005
R3674 VPWR.n1106 VPWR.n62 9.3005
R3675 VPWR.n1105 VPWR.n1104 9.3005
R3676 VPWR.n1103 VPWR.n63 9.3005
R3677 VPWR.n1103 VPWR.n64 9.3005
R3678 VPWR.n1102 VPWR.n67 9.3005
R3679 VPWR.n1101 VPWR.n68 9.3005
R3680 VPWR.n1100 VPWR.n1099 9.3005
R3681 VPWR.n1098 VPWR.n70 9.3005
R3682 VPWR.n1097 VPWR.n1096 9.3005
R3683 VPWR.n1095 VPWR.n72 9.3005
R3684 VPWR.n1094 VPWR.n73 9.3005
R3685 VPWR.n1093 VPWR.n1092 9.3005
R3686 VPWR.n1091 VPWR.n76 9.3005
R3687 VPWR.n1090 VPWR.n1089 9.3005
R3688 VPWR.n1088 VPWR.n1078 9.3005
R3689 VPWR.n910 VPWR.n909 9.3005
R3690 VPWR.n921 VPWR.n920 9.3005
R3691 VPWR.n925 VPWR.n924 9.3005
R3692 VPWR.n927 VPWR.n926 9.3005
R3693 VPWR.n928 VPWR.n330 9.3005
R3694 VPWR.n931 VPWR.n930 9.3005
R3695 VPWR.n932 VPWR.n329 9.3005
R3696 VPWR.n934 VPWR.n933 9.3005
R3697 VPWR.n935 VPWR.n328 9.3005
R3698 VPWR.n937 VPWR.n936 9.3005
R3699 VPWR.n939 VPWR.n938 9.3005
R3700 VPWR.n940 VPWR.n326 9.3005
R3701 VPWR.n943 VPWR.n942 9.3005
R3702 VPWR.n945 VPWR.n944 9.3005
R3703 VPWR.n948 VPWR.n947 9.3005
R3704 VPWR.n960 VPWR.n959 9.3005
R3705 VPWR.n961 VPWR.n317 9.3005
R3706 VPWR.n964 VPWR.n963 9.3005
R3707 VPWR.n965 VPWR.n316 9.3005
R3708 VPWR.n967 VPWR.n966 9.3005
R3709 VPWR.n968 VPWR.n315 9.3005
R3710 VPWR.n970 VPWR.n969 9.3005
R3711 VPWR.n972 VPWR.n971 9.3005
R3712 VPWR.n973 VPWR.n313 9.3005
R3713 VPWR.n976 VPWR.n975 9.3005
R3714 VPWR.n978 VPWR.n977 9.3005
R3715 VPWR.n980 VPWR.n979 9.3005
R3716 VPWR.n982 VPWR.n981 9.3005
R3717 VPWR.n983 VPWR.n309 9.3005
R3718 VPWR.n986 VPWR.n985 9.3005
R3719 VPWR.n990 VPWR.n97 9.3005
R3720 VPWR.n1001 VPWR.n1000 9.3005
R3721 VPWR.n1002 VPWR.n96 9.3005
R3722 VPWR.n1005 VPWR.n1004 9.3005
R3723 VPWR.n1007 VPWR.n1006 9.3005
R3724 VPWR.n1010 VPWR.n1009 9.3005
R3725 VPWR.n1011 VPWR.n94 9.3005
R3726 VPWR.n1013 VPWR.n1012 9.3005
R3727 VPWR.n1016 VPWR.n1015 9.3005
R3728 VPWR.n1018 VPWR.n1017 9.3005
R3729 VPWR.n1019 VPWR.n90 9.3005
R3730 VPWR.n1021 VPWR.n1020 9.3005
R3731 VPWR.n1023 VPWR.n1022 9.3005
R3732 VPWR.n1024 VPWR.n87 9.3005
R3733 VPWR.n1028 VPWR.n1027 9.3005
R3734 VPWR.n1030 VPWR.n1029 9.3005
R3735 VPWR.n1060 VPWR.n1059 9.3005
R3736 VPWR.n1058 VPWR.n1031 9.3005
R3737 VPWR.n1057 VPWR.n1056 9.3005
R3738 VPWR.n883 VPWR.n882 9.3005
R3739 VPWR.n698 VPWR.n432 9.3005
R3740 VPWR.n706 VPWR.n705 9.3005
R3741 VPWR.n708 VPWR.n707 9.3005
R3742 VPWR.n711 VPWR.n710 9.3005
R3743 VPWR.n713 VPWR.n712 9.3005
R3744 VPWR.n714 VPWR.n694 9.3005
R3745 VPWR.n717 VPWR.n716 9.3005
R3746 VPWR.n719 VPWR.n718 9.3005
R3747 VPWR.n720 VPWR.n692 9.3005
R3748 VPWR.n722 VPWR.n721 9.3005
R3749 VPWR.n723 VPWR.n691 9.3005
R3750 VPWR.n725 VPWR.n724 9.3005
R3751 VPWR.n726 VPWR.n690 9.3005
R3752 VPWR.n729 VPWR.n728 9.3005
R3753 VPWR.n731 VPWR.n730 9.3005
R3754 VPWR.n734 VPWR.n733 9.3005
R3755 VPWR.n745 VPWR.n744 9.3005
R3756 VPWR.n746 VPWR.n438 9.3005
R3757 VPWR.n749 VPWR.n748 9.3005
R3758 VPWR.n751 VPWR.n750 9.3005
R3759 VPWR.n752 VPWR.n436 9.3005
R3760 VPWR.n754 VPWR.n753 9.3005
R3761 VPWR.n755 VPWR.n435 9.3005
R3762 VPWR.n757 VPWR.n756 9.3005
R3763 VPWR.n758 VPWR.n434 9.3005
R3764 VPWR.n762 VPWR.n761 9.3005
R3765 VPWR.n763 VPWR.n433 9.3005
R3766 VPWR.n879 VPWR.n764 9.3005
R3767 VPWR.n878 VPWR.n766 9.3005
R3768 VPWR.n877 VPWR 9.3005
R3769 VPWR.n876 VPWR.n875 9.3005
R3770 VPWR.n775 VPWR.n772 9.3005
R3771 VPWR VPWR.n867 9.3005
R3772 VPWR.n866 VPWR.n865 9.3005
R3773 VPWR.n864 VPWR.n778 9.3005
R3774 VPWR.n863 VPWR.n862 9.3005
R3775 VPWR.n787 VPWR.n785 9.3005
R3776 VPWR.n857 VPWR 9.3005
R3777 VPWR.n856 VPWR.n790 9.3005
R3778 VPWR.n855 VPWR.n854 9.3005
R3779 VPWR.n852 VPWR.n851 9.3005
R3780 VPWR.n850 VPWR.n793 9.3005
R3781 VPWR.n849 VPWR.n848 9.3005
R3782 VPWR.n847 VPWR.n794 9.3005
R3783 VPWR.n845 VPWR.n844 9.3005
R3784 VPWR.n843 VPWR.n796 9.3005
R3785 VPWR.n842 VPWR.n841 9.3005
R3786 VPWR.n839 VPWR.n838 9.3005
R3787 VPWR.n810 VPWR.n802 9.3005
R3788 VPWR.n830 VPWR.n829 9.3005
R3789 VPWR.n828 VPWR.n827 9.3005
R3790 VPWR.n826 VPWR.n814 9.3005
R3791 VPWR.n825 VPWR.n824 9.3005
R3792 VPWR.n472 VPWR.n471 9.3005
R3793 VPWR.n475 VPWR.n461 9.3005
R3794 VPWR.n477 VPWR.n476 9.3005
R3795 VPWR.n547 VPWR.n546 9.3005
R3796 VPWR.n548 VPWR.n459 9.3005
R3797 VPWR.n484 VPWR.n458 9.3005
R3798 VPWR.n537 VPWR.n536 9.3005
R3799 VPWR.n534 VPWR.n486 9.3005
R3800 VPWR.n532 VPWR.n531 9.3005
R3801 VPWR.n530 VPWR.n491 9.3005
R3802 VPWR.n529 VPWR.n528 9.3005
R3803 VPWR.n526 VPWR.n492 9.3005
R3804 VPWR.n524 VPWR.n523 9.3005
R3805 VPWR.n522 VPWR.n521 9.3005
R3806 VPWR.n519 VPWR.n494 9.3005
R3807 VPWR.n518 VPWR.n517 9.3005
R3808 VPWR.n516 VPWR.n515 9.3005
R3809 VPWR.n513 VPWR.n496 9.3005
R3810 VPWR.n512 VPWR.n511 9.3005
R3811 VPWR.n510 VPWR.n497 9.3005
R3812 VPWR.n501 VPWR.n500 9.3005
R3813 VPWR.n502 VPWR.n450 9.3005
R3814 VPWR.n680 VPWR.n679 9.3005
R3815 VPWR.n677 VPWR.n449 9.3005
R3816 VPWR.n675 VPWR.n674 9.3005
R3817 VPWR.n673 VPWR.n672 9.3005
R3818 VPWR.n671 VPWR.n670 9.3005
R3819 VPWR.n669 VPWR.n453 9.3005
R3820 VPWR.n668 VPWR.n667 9.3005
R3821 VPWR.n666 VPWR.n454 9.3005
R3822 VPWR.n664 VPWR.n663 9.3005
R3823 VPWR.n662 VPWR.n457 9.3005
R3824 VPWR.n661 VPWR.n660 9.3005
R3825 VPWR.n659 VPWR.n658 9.3005
R3826 VPWR.n657 VPWR.n551 9.3005
R3827 VPWR.n656 VPWR.n655 9.3005
R3828 VPWR.n567 VPWR.n554 9.3005
R3829 VPWR.n563 VPWR.n556 9.3005
R3830 VPWR.n650 VPWR.n649 9.3005
R3831 VPWR.n648 VPWR.n557 9.3005
R3832 VPWR.n647 VPWR.n646 9.3005
R3833 VPWR.n645 VPWR.n576 9.3005
R3834 VPWR.n643 VPWR.n642 9.3005
R3835 VPWR.n641 VPWR.n578 9.3005
R3836 VPWR.n640 VPWR.n639 9.3005
R3837 VPWR.n638 VPWR.n579 9.3005
R3838 VPWR.n637 VPWR.n636 9.3005
R3839 VPWR.n635 VPWR.n634 9.3005
R3840 VPWR.n633 VPWR.n583 9.3005
R3841 VPWR.n632 VPWR.n631 9.3005
R3842 VPWR.n630 VPWR.n586 9.3005
R3843 VPWR.n629 VPWR.n628 9.3005
R3844 VPWR.n627 VPWR.n626 9.3005
R3845 VPWR.n592 VPWR.n590 9.3005
R3846 VPWR.n618 VPWR.n617 9.3005
R3847 VPWR.n616 VPWR.n601 9.3005
R3848 VPWR.n615 VPWR.n614 9.3005
R3849 VPWR.n613 VPWR.n604 9.3005
R3850 VPWR.n164 VPWR.n163 9.3005
R3851 VPWR.n166 VPWR.n165 9.3005
R3852 VPWR.n167 VPWR.n150 9.3005
R3853 VPWR.n171 VPWR.n170 9.3005
R3854 VPWR.n178 VPWR.n177 9.3005
R3855 VPWR.n6 VPWR.n0 9.3005
R3856 VPWR.n1191 VPWR.n1190 9.3005
R3857 VPWR.n1189 VPWR.n1188 9.3005
R3858 VPWR.n1187 VPWR.n1186 9.3005
R3859 VPWR.n1184 VPWR.n9 9.3005
R3860 VPWR.n1183 VPWR.n1182 9.3005
R3861 VPWR.n1181 VPWR.n1180 9.3005
R3862 VPWR.n1178 VPWR.n13 9.3005
R3863 VPWR.n1177 VPWR.n1176 9.3005
R3864 VPWR.n1175 VPWR.n1174 9.3005
R3865 VPWR.n1172 VPWR.n16 9.3005
R3866 VPWR.n1171 VPWR.n1170 9.3005
R3867 VPWR.n1169 VPWR.n18 9.3005
R3868 VPWR.n1168 VPWR.n1167 9.3005
R3869 VPWR.n1166 VPWR.n1165 9.3005
R3870 VPWR.n125 VPWR.n22 9.3005
R3871 VPWR.n135 VPWR.n134 9.3005
R3872 VPWR.n137 VPWR.n136 9.3005
R3873 VPWR.n140 VPWR.n139 9.3005
R3874 VPWR.n141 VPWR.n115 9.3005
R3875 VPWR.n142 VPWR.n112 9.3005
R3876 VPWR.n143 VPWR.n111 9.3005
R3877 VPWR.n145 VPWR.n144 9.3005
R3878 VPWR.n146 VPWR.n109 9.3005
R3879 VPWR.n181 VPWR.n147 9.3005
R3880 VPWR.n183 VPWR.n182 9.3005
R3881 VPWR.n184 VPWR.n108 9.3005
R3882 VPWR.n187 VPWR.n185 9.3005
R3883 VPWR.n285 VPWR.n284 9.3005
R3884 VPWR.n283 VPWR.n189 9.3005
R3885 VPWR.n282 VPWR.n197 9.3005
R3886 VPWR.n281 VPWR.n200 9.3005
R3887 VPWR.n280 VPWR.n279 9.3005
R3888 VPWR.n278 VPWR.n277 9.3005
R3889 VPWR.n275 VPWR.n274 9.3005
R3890 VPWR.n273 VPWR.n272 9.3005
R3891 VPWR.n270 VPWR.n205 9.3005
R3892 VPWR.n267 VPWR.n266 9.3005
R3893 VPWR.n265 VPWR.n208 9.3005
R3894 VPWR.n264 VPWR.n263 9.3005
R3895 VPWR.n261 VPWR.n260 9.3005
R3896 VPWR.n259 VPWR.n213 9.3005
R3897 VPWR.n258 VPWR.n257 9.3005
R3898 VPWR.n256 VPWR.n214 9.3005
R3899 VPWR.n255 VPWR.n254 9.3005
R3900 VPWR.n219 VPWR.n217 9.3005
R3901 VPWR.n246 VPWR.n245 9.3005
R3902 VPWR.n244 VPWR.n229 9.3005
R3903 VPWR.n243 VPWR.n242 9.3005
R3904 VPWR.n241 VPWR.n232 9.3005
R3905 VPWR.n380 VPWR.n367 9.09802
R3906 VPWR.n1140 VPWR.n39 9.09802
R3907 VPWR.n1015 VPWR.n92 9.09802
R3908 VPWR.n1186 VPWR.n10 9.09802
R3909 VPWR.n1186 VPWR.n1185 9.09802
R3910 VPWR.n1174 VPWR.n1173 9.09802
R3911 VPWR.n879 VPWR.n433 9.03579
R3912 VPWR.n654 VPWR.n653 8.9761
R3913 VPWR.n1179 VPWR.n1178 8.56909
R3914 VPWR.n979 VPWR.n978 8.44958
R3915 VPWR.t415 VPWR.t443 8.39273
R3916 VPWR.t222 VPWR.t396 8.39273
R3917 VPWR.t337 VPWR.t104 8.39273
R3918 VPWR.t314 VPWR.t251 8.39273
R3919 VPWR.t427 VPWR.t464 8.39273
R3920 VPWR.t0 VPWR.t458 8.39273
R3921 VPWR.t94 VPWR.t345 8.39273
R3922 VPWR.n142 VPWR.n141 8.28285
R3923 VPWR.n135 VPWR.n22 8.28285
R3924 VPWR.n283 VPWR.n282 8.28285
R3925 VPWR.n357 VPWR.n342 7.98741
R3926 VPWR VPWR.n637 7.93438
R3927 VPWR.n582 VPWR.n581 7.93438
R3928 VPWR.n20 VPWR.n19 7.93438
R3929 VPWR.n983 VPWR.n982 7.75995
R3930 VPWR.n643 VPWR.n578 7.75995
R3931 VPWR.n940 VPWR.n939 7.21067
R3932 VPWR.n947 VPWR.n945 7.21067
R3933 VPWR.n973 VPWR.n972 7.21067
R3934 VPWR.n1114 VPWR.n56 7.11161
R3935 VPWR.n846 VPWR.n845 7.0168
R3936 VPWR.n705 VPWR.n696 6.85159
R3937 VPWR.t32 VPWR.t389 6.71428
R3938 VPWR.t357 VPWR.t8 6.71428
R3939 VPWR.n405 VPWR.n358 6.66496
R3940 VPWR.n1142 VPWR.n1141 6.66496
R3941 VPWR.n1009 VPWR.n1008 6.66496
R3942 VPWR.n672 VPWR.n451 6.66496
R3943 VPWR.n553 VPWR.n551 6.66496
R3944 VPWR.n1020 VPWR.n89 6.45339
R3945 VPWR.n380 VPWR.n379 6.34761
R3946 VPWR.n1153 VPWR.n36 6.34761
R3947 VPWR.n526 VPWR.n525 6.16836
R3948 VPWR.n1027 VPWR.n1026 6.13604
R3949 VPWR.n760 VPWR.n433 6.12224
R3950 VPWR.n928 VPWR.n927 5.66204
R3951 VPWR.n930 VPWR.n928 5.66204
R3952 VPWR.n934 VPWR.n329 5.66204
R3953 VPWR.n935 VPWR.n934 5.66204
R3954 VPWR.n936 VPWR.n935 5.66204
R3955 VPWR.n961 VPWR.n960 5.66204
R3956 VPWR.n963 VPWR.n961 5.66204
R3957 VPWR.n967 VPWR.n316 5.66204
R3958 VPWR.n968 VPWR.n967 5.66204
R3959 VPWR.n969 VPWR.n968 5.66204
R3960 VPWR.n746 VPWR.n745 5.66204
R3961 VPWR.n752 VPWR.n751 5.66204
R3962 VPWR.n753 VPWR.n752 5.66204
R3963 VPWR.n753 VPWR.n435 5.66204
R3964 VPWR.n757 VPWR.n435 5.66204
R3965 VPWR.n758 VPWR.n757 5.66204
R3966 VPWR.n714 VPWR.n713 5.66204
R3967 VPWR.n720 VPWR.n719 5.66204
R3968 VPWR.n721 VPWR.n720 5.66204
R3969 VPWR.n721 VPWR.n691 5.66204
R3970 VPWR.n725 VPWR.n691 5.66204
R3971 VPWR.n726 VPWR.n725 5.66204
R3972 VPWR.n519 VPWR.n518 5.66204
R3973 VPWR.n513 VPWR.n512 5.66204
R3974 VPWR.n512 VPWR.n497 5.66204
R3975 VPWR.n500 VPWR.n497 5.66204
R3976 VPWR.n500 VPWR.n450 5.66204
R3977 VPWR.n679 VPWR.n450 5.66204
R3978 VPWR.n728 VPWR.n689 5.48759
R3979 VPWR.n677 VPWR.n676 5.48759
R3980 VPWR.n924 VPWR.n922 5.42606
R3981 VPWR.n733 VPWR.n732 5.42606
R3982 VPWR.n710 VPWR.n709 5.42606
R3983 VPWR.n521 VPWR.n493 5.42606
R3984 VPWR.n902 VPWR.n901 5.40233
R3985 VPWR.n425 VPWR.n424 5.40233
R3986 VPWR.n665 VPWR.n456 5.40233
R3987 VPWR.n936 VPWR.n327 5.29281
R3988 VPWR.n942 VPWR.n941 5.29281
R3989 VPWR.n942 VPWR.n325 5.29281
R3990 VPWR.n969 VPWR.n314 5.29281
R3991 VPWR.n975 VPWR.n974 5.29281
R3992 VPWR.n975 VPWR.n312 5.29281
R3993 VPWR.n745 VPWR.n439 5.29281
R3994 VPWR.n759 VPWR.n758 5.29281
R3995 VPWR.n713 VPWR.n695 5.29281
R3996 VPWR.n727 VPWR.n726 5.29281
R3997 VPWR.n520 VPWR.n519 5.29281
R3998 VPWR.n679 VPWR.n678 5.29281
R3999 VPWR.n346 VPWR.n345 5.25888
R4000 VPWR.n377 VPWR.n370 5.18397
R4001 VPWR.n979 VPWR.n310 5.18397
R4002 VPWR.n1014 VPWR.n1013 5.18397
R4003 VPWR.n455 VPWR.n453 5.18397
R4004 VPWR.n1183 VPWR.n12 5.18397
R4005 VPWR.t13 VPWR.t417 5.03584
R4006 VPWR.t277 VPWR.t462 5.03584
R4007 VPWR.t4 VPWR.t305 5.03584
R4008 VPWR.t399 VPWR.t343 5.03584
R4009 VPWR.t285 VPWR.t355 5.03584
R4010 VPWR.n652 VPWR.n651 5.00648
R4011 VPWR.n404 VPWR.n359 4.98946
R4012 VPWR.n921 VPWR.n333 4.94058
R4013 VPWR.n533 VPWR.n490 4.92694
R4014 VPWR.n666 VPWR.n665 4.86662
R4015 VPWR.n665 VPWR.n664 4.86662
R4016 VPWR.n1004 VPWR.n95 4.79796
R4017 VPWR.n344 VPWR.n343 4.77455
R4018 VPWR.n1132 VPWR.n1131 4.67352
R4019 VPWR.n882 VPWR.n432 4.67352
R4020 VPWR.n705 VPWR.n432 4.67352
R4021 VPWR.n867 VPWR.n866 4.67352
R4022 VPWR.n866 VPWR.n778 4.67352
R4023 VPWR.n829 VPWR.n810 4.67352
R4024 VPWR.n829 VPWR.n828 4.67352
R4025 VPWR.n828 VPWR.n814 4.67352
R4026 VPWR.n476 VPWR.n475 4.67352
R4027 VPWR.n167 VPWR.n166 4.67352
R4028 VPWR.n355 VPWR.n346 4.62124
R4029 VPWR.n357 VPWR.n356 4.62124
R4030 VPWR.n921 VPWR.n332 4.62124
R4031 VPWR.n488 VPWR.n487 4.5918
R4032 VPWR.n982 VPWR.n310 4.54926
R4033 VPWR.n1015 VPWR.n1014 4.54926
R4034 VPWR.n667 VPWR.n455 4.54926
R4035 VPWR.n1180 VPWR.n12 4.54926
R4036 VPWR.n174 VPWR.n172 4.51401
R4037 VPWR.n1193 VPWR.n1192 4.51401
R4038 VPWR.n1164 VPWR.n1163 4.51401
R4039 VPWR.n131 VPWR.n122 4.51401
R4040 VPWR.n288 VPWR.n105 4.51401
R4041 VPWR.n196 VPWR.n195 4.51401
R4042 VPWR.n1158 VPWR.n31 4.51401
R4043 VPWR.n1149 VPWR.n1145 4.51401
R4044 VPWR.n409 VPWR.n339 4.51401
R4045 VPWR.n400 VPWR.n399 4.51401
R4046 VPWR.n1072 VPWR.n71 4.51401
R4047 VPWR.n1077 VPWR.n1076 4.51401
R4048 VPWR.n304 VPWR.n293 4.51401
R4049 VPWR.n294 VPWR.n57 4.51401
R4050 VPWR.n951 VPWR.n324 4.51401
R4051 VPWR.n956 VPWR.n320 4.51401
R4052 VPWR.n913 VPWR.n890 4.51401
R4053 VPWR.n917 VPWR.n334 4.51401
R4054 VPWR.n1063 VPWR.n84 4.51401
R4055 VPWR.n1046 VPWR.n1045 4.51401
R4056 VPWR.n993 VPWR.n987 4.51401
R4057 VPWR.n997 VPWR.n99 4.51401
R4058 VPWR.n570 VPWR.n552 4.51401
R4059 VPWR.n575 VPWR.n574 4.51401
R4060 VPWR.n874 VPWR.n873 4.51401
R4061 VPWR.n784 VPWR.n783 4.51401
R4062 VPWR.n886 VPWR.n415 4.51401
R4063 VPWR.n704 VPWR.n703 4.51401
R4064 VPWR.n806 VPWR.n797 4.51401
R4065 VPWR.n832 VPWR.n831 4.51401
R4066 VPWR.n737 VPWR.n686 4.51401
R4067 VPWR.n741 VPWR.n441 4.51401
R4068 VPWR.n509 VPWR.n508 4.51401
R4069 VPWR.n682 VPWR.n681 4.51401
R4070 VPWR.n597 VPWR.n587 4.51401
R4071 VPWR.n620 VPWR.n619 4.51401
R4072 VPWR.n545 VPWR.n544 4.51401
R4073 VPWR.n539 VPWR.n538 4.51401
R4074 VPWR.n224 VPWR.n222 4.51401
R4075 VPWR.n248 VPWR.n247 4.51401
R4076 VPWR.n408 VPWR.n407 4.5005
R4077 VPWR.n360 VPWR 4.5005
R4078 VPWR.n402 VPWR.n401 4.5005
R4079 VPWR.n1157 VPWR.n1156 4.5005
R4080 VPWR.n1146 VPWR.n33 4.5005
R4081 VPWR.n1151 VPWR.n1150 4.5005
R4082 VPWR.n1071 VPWR.n1070 4.5005
R4083 VPWR.n1068 VPWR 4.5005
R4084 VPWR.n78 VPWR.n77 4.5005
R4085 VPWR.n303 VPWR.n302 4.5005
R4086 VPWR.n300 VPWR.n299 4.5005
R4087 VPWR.n296 VPWR.n295 4.5005
R4088 VPWR.n912 VPWR.n911 4.5005
R4089 VPWR.n891 VPWR 4.5005
R4090 VPWR.n919 VPWR.n918 4.5005
R4091 VPWR.n950 VPWR.n949 4.5005
R4092 VPWR.n322 VPWR.n319 4.5005
R4093 VPWR.n958 VPWR.n957 4.5005
R4094 VPWR.n1062 VPWR.n1061 4.5005
R4095 VPWR.n1041 VPWR.n1040 4.5005
R4096 VPWR.n1044 VPWR.n1039 4.5005
R4097 VPWR.n992 VPWR.n991 4.5005
R4098 VPWR.n988 VPWR.n98 4.5005
R4099 VPWR.n999 VPWR.n998 4.5005
R4100 VPWR.n885 VPWR.n884 4.5005
R4101 VPWR.n699 VPWR 4.5005
R4102 VPWR.n702 VPWR.n697 4.5005
R4103 VPWR.n771 VPWR.n768 4.5005
R4104 VPWR.n869 VPWR.n868 4.5005
R4105 VPWR.n780 VPWR.n779 4.5005
R4106 VPWR.n805 VPWR.n801 4.5005
R4107 VPWR.n837 VPWR.n836 4.5005
R4108 VPWR.n809 VPWR.n804 4.5005
R4109 VPWR.n736 VPWR.n735 4.5005
R4110 VPWR.n687 VPWR.n440 4.5005
R4111 VPWR.n743 VPWR.n742 4.5005
R4112 VPWR.n507 VPWR.n498 4.5005
R4113 VPWR.n504 VPWR.n503 4.5005
R4114 VPWR.n448 VPWR.n447 4.5005
R4115 VPWR.n569 VPWR.n568 4.5005
R4116 VPWR.n566 VPWR.n565 4.5005
R4117 VPWR.n559 VPWR.n558 4.5005
R4118 VPWR.n596 VPWR.n591 4.5005
R4119 VPWR.n625 VPWR.n624 4.5005
R4120 VPWR.n600 VPWR.n594 4.5005
R4121 VPWR.n479 VPWR.n478 4.5005
R4122 VPWR VPWR.n483 4.5005
R4123 VPWR.n485 VPWR.n482 4.5005
R4124 VPWR.n176 VPWR.n175 4.5005
R4125 VPWR VPWR.n1197 4.5005
R4126 VPWR.n5 VPWR.n2 4.5005
R4127 VPWR.n124 VPWR.n24 4.5005
R4128 VPWR.n128 VPWR.n126 4.5005
R4129 VPWR.n133 VPWR.n132 4.5005
R4130 VPWR.n287 VPWR.n286 4.5005
R4131 VPWR.n191 VPWR 4.5005
R4132 VPWR.n194 VPWR.n190 4.5005
R4133 VPWR.n223 VPWR.n218 4.5005
R4134 VPWR.n253 VPWR.n252 4.5005
R4135 VPWR.n228 VPWR.n221 4.5005
R4136 VPWR.n1119 VPWR.n1118 4.36875
R4137 VPWR.n867 VPWR.n777 4.36875
R4138 VPWR.n862 VPWR.n786 4.36875
R4139 VPWR.n862 VPWR.n861 4.36875
R4140 VPWR.n810 VPWR.n800 4.36875
R4141 VPWR.n815 VPWR.n814 4.36875
R4142 VPWR.n476 VPWR.n460 4.36875
R4143 VPWR.n169 VPWR.n168 4.26717
R4144 VPWR.n353 VPWR.n349 4.02033
R4145 VPWR.n353 VPWR.n352 4.02033
R4146 VPWR.n1087 VPWR.n1082 4.02033
R4147 VPWR.n1087 VPWR.n1085 4.02033
R4148 VPWR.n900 VPWR.n896 4.02033
R4149 VPWR.n900 VPWR.n899 4.02033
R4150 VPWR.n1038 VPWR.n1035 4.02033
R4151 VPWR.n1053 VPWR.n1049 4.02033
R4152 VPWR.n1053 VPWR.n1052 4.02033
R4153 VPWR.n423 VPWR.n419 4.02033
R4154 VPWR.n423 VPWR.n422 4.02033
R4155 VPWR.n823 VPWR.n818 4.02033
R4156 VPWR.n823 VPWR.n821 4.02033
R4157 VPWR.n469 VPWR.n465 4.02033
R4158 VPWR.n469 VPWR.n468 4.02033
R4159 VPWR.n611 VPWR.n607 4.02033
R4160 VPWR.n611 VPWR.n610 4.02033
R4161 VPWR.n121 VPWR.n118 4.02033
R4162 VPWR.n160 VPWR.n155 4.02033
R4163 VPWR.n160 VPWR.n159 4.02033
R4164 VPWR.n239 VPWR.n235 4.02033
R4165 VPWR.n239 VPWR.n238 4.02033
R4166 VPWR.n358 VPWR.n357 3.78037
R4167 VPWR.n277 VPWR.n201 3.76521
R4168 VPWR.n263 VPWR.n209 3.76521
R4169 VPWR.n1119 VPWR.n52 3.50526
R4170 VPWR.n393 VPWR.n364 3.47425
R4171 VPWR.n389 VPWR.n364 3.47425
R4172 VPWR.n389 VPWR.n388 3.47425
R4173 VPWR.n388 VPWR.n387 3.47425
R4174 VPWR.n985 VPWR.n97 3.47425
R4175 VPWR.n1001 VPWR.n97 3.47425
R4176 VPWR.n1002 VPWR.n1001 3.47425
R4177 VPWR.n650 VPWR.n557 3.47425
R4178 VPWR.n646 VPWR.n645 3.47425
R4179 VPWR.n1194 VPWR.n1193 3.43925
R4180 VPWR.n174 VPWR.n173 3.43925
R4181 VPWR.n131 VPWR.n27 3.43925
R4182 VPWR.n1163 VPWR.n1162 3.43925
R4183 VPWR.n195 VPWR.n103 3.43925
R4184 VPWR.n289 VPWR.n288 3.43925
R4185 VPWR.n1149 VPWR.n28 3.43925
R4186 VPWR.n1159 VPWR.n1158 3.43925
R4187 VPWR.n400 VPWR.n337 3.43925
R4188 VPWR.n410 VPWR.n409 3.43925
R4189 VPWR.n1076 VPWR.n1075 3.43925
R4190 VPWR.n1073 VPWR.n1072 3.43925
R4191 VPWR.n294 VPWR.n291 3.43925
R4192 VPWR.n305 VPWR.n304 3.43925
R4193 VPWR.n956 VPWR.n955 3.43925
R4194 VPWR.n952 VPWR.n951 3.43925
R4195 VPWR.n917 VPWR.n916 3.43925
R4196 VPWR.n914 VPWR.n913 3.43925
R4197 VPWR.n1045 VPWR.n81 3.43925
R4198 VPWR.n1064 VPWR.n1063 3.43925
R4199 VPWR.n997 VPWR.n996 3.43925
R4200 VPWR.n994 VPWR.n993 3.43925
R4201 VPWR.n574 VPWR.n573 3.43925
R4202 VPWR.n571 VPWR.n570 3.43925
R4203 VPWR.n703 VPWR.n412 3.43925
R4204 VPWR.n887 VPWR.n886 3.43925
R4205 VPWR.n833 VPWR.n832 3.43925
R4206 VPWR.n807 VPWR.n806 3.43925
R4207 VPWR.n741 VPWR.n740 3.43925
R4208 VPWR.n738 VPWR.n737 3.43925
R4209 VPWR.n621 VPWR.n620 3.43925
R4210 VPWR.n598 VPWR.n597 3.43925
R4211 VPWR.n540 VPWR.n539 3.43925
R4212 VPWR.n544 VPWR.n543 3.43925
R4213 VPWR.n3 VPWR.n1 3.4105
R4214 VPWR.n1196 VPWR.n1195 3.4105
R4215 VPWR.n127 VPWR.n25 3.4105
R4216 VPWR.n130 VPWR.n129 3.4105
R4217 VPWR.n106 VPWR.n104 3.4105
R4218 VPWR.n193 VPWR.n192 3.4105
R4219 VPWR.n32 VPWR.n30 3.4105
R4220 VPWR.n1148 VPWR.n1147 3.4105
R4221 VPWR.n340 VPWR.n338 3.4105
R4222 VPWR.n362 VPWR.n361 3.4105
R4223 VPWR.n1069 VPWR.n1066 3.4105
R4224 VPWR.n1067 VPWR.n79 3.4105
R4225 VPWR.n301 VPWR.n292 3.4105
R4226 VPWR.n298 VPWR.n297 3.4105
R4227 VPWR.n953 VPWR.n323 3.4105
R4228 VPWR.n954 VPWR.n321 3.4105
R4229 VPWR.n892 VPWR.n889 3.4105
R4230 VPWR.n336 VPWR.n335 3.4105
R4231 VPWR.n85 VPWR.n83 3.4105
R4232 VPWR.n1043 VPWR.n1042 3.4105
R4233 VPWR.n989 VPWR.n308 3.4105
R4234 VPWR.n101 VPWR.n100 3.4105
R4235 VPWR.n562 VPWR.n561 3.4105
R4236 VPWR.n564 VPWR.n560 3.4105
R4237 VPWR.n782 VPWR.n307 3.4105
R4238 VPWR.n872 VPWR.n307 3.4105
R4239 VPWR.n783 VPWR.n782 3.4105
R4240 VPWR.n873 VPWR.n872 3.4105
R4241 VPWR.n871 VPWR.n870 3.4105
R4242 VPWR.n781 VPWR.n770 3.4105
R4243 VPWR.n416 VPWR.n414 3.4105
R4244 VPWR.n701 VPWR.n700 3.4105
R4245 VPWR.n808 VPWR.n803 3.4105
R4246 VPWR.n835 VPWR.n834 3.4105
R4247 VPWR.n688 VPWR.n685 3.4105
R4248 VPWR.n443 VPWR.n442 3.4105
R4249 VPWR.n684 VPWR.n683 3.4105
R4250 VPWR.n684 VPWR.n445 3.4105
R4251 VPWR.n683 VPWR.n682 3.4105
R4252 VPWR.n508 VPWR.n445 3.4105
R4253 VPWR.n506 VPWR.n505 3.4105
R4254 VPWR.n499 VPWR.n446 3.4105
R4255 VPWR.n595 VPWR.n593 3.4105
R4256 VPWR.n623 VPWR.n622 3.4105
R4257 VPWR.n542 VPWR.n480 3.4105
R4258 VPWR.n541 VPWR.n481 3.4105
R4259 VPWR.n249 VPWR.n80 3.4105
R4260 VPWR.n225 VPWR.n80 3.4105
R4261 VPWR.n249 VPWR.n248 3.4105
R4262 VPWR.n225 VPWR.n224 3.4105
R4263 VPWR.n226 VPWR.n220 3.4105
R4264 VPWR.n251 VPWR.n250 3.4105
R4265 VPWR.n269 VPWR.n268 3.38874
R4266 VPWR.n379 VPWR.n378 3.38562
R4267 VPWR.n1143 VPWR.n36 3.38562
R4268 VPWR.n651 VPWR.n650 3.36097
R4269 VPWR.t241 VPWR.t411 3.35739
R4270 VPWR.t259 VPWR.t351 3.35739
R4271 VPWR.n1023 VPWR.n89 3.27984
R4272 VPWR.n396 VPWR.n395 3.2477
R4273 VPWR.n387 VPWR.n366 3.2477
R4274 VPWR.n985 VPWR.n984 3.2477
R4275 VPWR.n1003 VPWR.n1002 3.2477
R4276 VPWR.n556 VPWR.n555 3.2477
R4277 VPWR.n645 VPWR.n644 3.2477
R4278 VPWR.n1131 VPWR.n1130 3.2005
R4279 VPWR.n814 VPWR.n813 3.12116
R4280 VPWR.n374 VPWR.n373 3.06827
R4281 VPWR.n1141 VPWR.n1140 3.06827
R4282 VPWR.n354 VPWR.n353 3.05586
R4283 VPWR.n903 VPWR.n900 3.05586
R4284 VPWR.n426 VPWR.n423 3.05586
R4285 VPWR.n470 VPWR.n469 3.05586
R4286 VPWR.n160 VPWR.n156 3.05586
R4287 VPWR.n1087 VPWR.n1086 3.04861
R4288 VPWR.n1054 VPWR.n1053 3.04861
R4289 VPWR.n1055 VPWR.n1038 3.04861
R4290 VPWR.n823 VPWR.n822 3.04861
R4291 VPWR.n612 VPWR.n611 3.04861
R4292 VPWR.n240 VPWR.n239 3.04861
R4293 VPWR.n138 VPWR.n121 3.04861
R4294 VPWR.n930 VPWR.n929 3.01588
R4295 VPWR.n963 VPWR.n962 3.01588
R4296 VPWR.n747 VPWR.n746 3.01588
R4297 VPWR.n748 VPWR.n437 3.01588
R4298 VPWR.n715 VPWR.n714 3.01588
R4299 VPWR.n716 VPWR.n693 3.01588
R4300 VPWR.n518 VPWR.n495 3.01588
R4301 VPWR.n515 VPWR.n514 3.01588
R4302 VPWR.n882 VPWR.n431 2.99733
R4303 VPWR.n1026 VPWR.n86 2.96248
R4304 VPWR.n906 VPWR.n905 2.87861
R4305 VPWR.n429 VPWR.n428 2.87861
R4306 VPWR.n397 VPWR.n359 2.69393
R4307 VPWR.n923 VPWR.n331 2.64665
R4308 VPWR.n927 VPWR.n331 2.64665
R4309 VPWR.n929 VPWR.n329 2.64665
R4310 VPWR.n946 VPWR.n318 2.64665
R4311 VPWR.n960 VPWR.n318 2.64665
R4312 VPWR.n962 VPWR.n316 2.64665
R4313 VPWR.n748 VPWR.n747 2.64665
R4314 VPWR.n751 VPWR.n437 2.64665
R4315 VPWR.n716 VPWR.n715 2.64665
R4316 VPWR.n719 VPWR.n693 2.64665
R4317 VPWR.n515 VPWR.n495 2.64665
R4318 VPWR.n514 VPWR.n513 2.64665
R4319 VPWR.n813 VPWR.n811 2.63539
R4320 VPWR.n349 VPWR.n347 2.63539
R4321 VPWR.n352 VPWR.n350 2.63539
R4322 VPWR.n1082 VPWR.n1080 2.63539
R4323 VPWR.n1085 VPWR.n1083 2.63539
R4324 VPWR.n896 VPWR.n894 2.63539
R4325 VPWR.n899 VPWR.n897 2.63539
R4326 VPWR.n1035 VPWR.n1033 2.63539
R4327 VPWR.n1049 VPWR.n1047 2.63539
R4328 VPWR.n1052 VPWR.n1050 2.63539
R4329 VPWR.n419 VPWR.n417 2.63539
R4330 VPWR.n422 VPWR.n420 2.63539
R4331 VPWR.n818 VPWR.n816 2.63539
R4332 VPWR.n821 VPWR.n819 2.63539
R4333 VPWR.n465 VPWR.n463 2.63539
R4334 VPWR.n468 VPWR.n466 2.63539
R4335 VPWR.n607 VPWR.n605 2.63539
R4336 VPWR.n610 VPWR.n608 2.63539
R4337 VPWR.n118 VPWR.n116 2.63539
R4338 VPWR.n155 VPWR.n153 2.63539
R4339 VPWR.n159 VPWR.n157 2.63539
R4340 VPWR.n235 VPWR.n233 2.63539
R4341 VPWR.n238 VPWR.n236 2.63539
R4342 VPWR.n908 VPWR.n907 2.61352
R4343 VPWR.n431 VPWR.n430 2.61352
R4344 VPWR.n532 VPWR.n491 2.50603
R4345 VPWR.n528 VPWR.n491 2.50603
R4346 VPWR.n533 VPWR.n532 2.45156
R4347 VPWR.n812 VPWR.n811 2.37495
R4348 VPWR.n351 VPWR.n350 2.37495
R4349 VPWR.n348 VPWR.n347 2.37495
R4350 VPWR.n1084 VPWR.n1083 2.37495
R4351 VPWR.n1081 VPWR.n1080 2.37495
R4352 VPWR.n898 VPWR.n897 2.37495
R4353 VPWR.n895 VPWR.n894 2.37495
R4354 VPWR.n1034 VPWR.n1033 2.37495
R4355 VPWR.n1051 VPWR.n1050 2.37495
R4356 VPWR.n1048 VPWR.n1047 2.37495
R4357 VPWR.n421 VPWR.n420 2.37495
R4358 VPWR.n418 VPWR.n417 2.37495
R4359 VPWR.n820 VPWR.n819 2.37495
R4360 VPWR.n817 VPWR.n816 2.37495
R4361 VPWR.n467 VPWR.n466 2.37495
R4362 VPWR.n464 VPWR.n463 2.37495
R4363 VPWR.n609 VPWR.n608 2.37495
R4364 VPWR.n606 VPWR.n605 2.37495
R4365 VPWR.n117 VPWR.n116 2.37495
R4366 VPWR.n158 VPWR.n157 2.37495
R4367 VPWR.n154 VPWR.n153 2.37495
R4368 VPWR.n237 VPWR.n236 2.37495
R4369 VPWR.n234 VPWR.n233 2.37495
R4370 VPWR.n535 VPWR.n534 2.34263
R4371 VPWR.n528 VPWR.n527 2.34263
R4372 VPWR.n475 VPWR.n474 2.33701
R4373 VPWR.n166 VPWR.n152 2.33701
R4374 VPWR.n922 VPWR.n921 2.28432
R4375 VPWR.n345 VPWR.n343 2.28374
R4376 VPWR.n178 VPWR.n149 2.25932
R4377 VPWR.n277 VPWR.n276 2.25932
R4378 VPWR.n272 VPWR.n271 2.25932
R4379 VPWR.n263 VPWR.n262 2.25932
R4380 VPWR.n905 VPWR.n904 2.25312
R4381 VPWR.n428 VPWR.n427 2.25312
R4382 VPWR.n44 VPWR.n43 2.03225
R4383 VPWR.n474 VPWR.n473 2.03225
R4384 VPWR.n577 VPWR.n557 1.85065
R4385 VPWR.n395 VPWR.n394 1.81289
R4386 VPWR.n638 VPWR 1.79885
R4387 VPWR.n761 VPWR.n760 1.78512
R4388 VPWR.n161 VPWR.n152 1.77828
R4389 VPWR.n847 VPWR.n846 1.70717
R4390 VPWR.n573 VPWR.n572 1.69188
R4391 VPWR.n572 VPWR.n571 1.69188
R4392 VPWR.n996 VPWR.n995 1.69188
R4393 VPWR.n995 VPWR.n994 1.69188
R4394 VPWR.n306 VPWR.n291 1.69188
R4395 VPWR.n306 VPWR.n305 1.69188
R4396 VPWR.n290 VPWR.n103 1.69188
R4397 VPWR.n290 VPWR.n289 1.69188
R4398 VPWR.n769 VPWR.n307 1.69188
R4399 VPWR.n740 VPWR.n739 1.69188
R4400 VPWR.n739 VPWR.n738 1.69188
R4401 VPWR.n955 VPWR.n29 1.69188
R4402 VPWR.n952 VPWR.n29 1.69188
R4403 VPWR.n1160 VPWR.n28 1.69188
R4404 VPWR.n1160 VPWR.n1159 1.69188
R4405 VPWR.n1161 VPWR.n27 1.69188
R4406 VPWR.n1162 VPWR.n1161 1.69188
R4407 VPWR.n684 VPWR.n444 1.69188
R4408 VPWR.n540 VPWR.n413 1.69188
R4409 VPWR.n543 VPWR.n413 1.69188
R4410 VPWR.n888 VPWR.n412 1.69188
R4411 VPWR.n888 VPWR.n887 1.69188
R4412 VPWR.n916 VPWR.n915 1.69188
R4413 VPWR.n915 VPWR.n914 1.69188
R4414 VPWR.n411 VPWR.n337 1.69188
R4415 VPWR.n411 VPWR.n410 1.69188
R4416 VPWR.n1194 VPWR.n4 1.69188
R4417 VPWR.n173 VPWR.n4 1.69188
R4418 VPWR.n621 VPWR.n599 1.69188
R4419 VPWR.n599 VPWR.n598 1.69188
R4420 VPWR.n833 VPWR.n82 1.69188
R4421 VPWR.n807 VPWR.n82 1.69188
R4422 VPWR.n1065 VPWR.n81 1.69188
R4423 VPWR.n1065 VPWR.n1064 1.69188
R4424 VPWR.n1075 VPWR.n1074 1.69188
R4425 VPWR.n1074 VPWR.n1073 1.69188
R4426 VPWR.n227 VPWR.n80 1.69188
R4427 VPWR VPWR.t474 1.67895
R4428 VPWR.t76 VPWR.t384 1.67895
R4429 VPWR.t283 VPWR.t84 1.67895
R4430 VPWR.n394 VPWR.n393 1.66186
R4431 VPWR.n1132 VPWR.n45 1.6259
R4432 VPWR.n646 VPWR.n577 1.6241
R4433 VPWR.n1111 VPWR.n56 1.61235
R4434 VPWR.n1124 VPWR.n1123 1.50638
R4435 VPWR.n373 VPWR.n370 1.48149
R4436 VPWR.n775 VPWR.n767 1.47352
R4437 VPWR.n858 VPWR.n787 1.47352
R4438 VPWR.n343 VPWR.n342 1.37322
R4439 VPWR.n908 VPWR.n906 1.2502
R4440 VPWR.n431 VPWR.n429 1.2502
R4441 VPWR.n1130 VPWR.n1129 1.16875
R4442 VPWR.n637 VPWR.n581 1.16414
R4443 VPWR.n1180 VPWR.n1179 1.16414
R4444 VPWR.n19 VPWR.n18 1.16414
R4445 VPWR.n841 VPWR.n840 1.12991
R4446 VPWR.n1038 VPWR.n1037 0.899674
R4447 VPWR.n121 VPWR.n120 0.899674
R4448 VPWR.n52 VPWR.n50 0.863992
R4449 VPWR.n908 VPWR.n333 0.848662
R4450 VPWR.n536 VPWR.n487 0.790287
R4451 VPWR.n45 VPWR.n44 0.711611
R4452 VPWR.n905 VPWR.n902 0.644287
R4453 VPWR.n428 VPWR.n425 0.644287
R4454 VPWR.n383 VPWR.n367 0.635211
R4455 VPWR.n1137 VPWR.n39 0.635211
R4456 VPWR.n1018 VPWR.n92 0.635211
R4457 VPWR.n1030 VPWR.n86 0.635211
R4458 VPWR.n634 VPWR.n582 0.635211
R4459 VPWR.n1185 VPWR.n1184 0.635211
R4460 VPWR.n1173 VPWR.n1172 0.635211
R4461 VPWR.n1167 VPWR.n20 0.635211
R4462 VPWR.n10 VPWR.n8 0.42364
R4463 VPWR.n853 VPWR.n852 0.376971
R4464 VPWR.n272 VPWR.n204 0.376971
R4465 VPWR.n268 VPWR.n267 0.376971
R4466 VPWR.n924 VPWR.n923 0.369731
R4467 VPWR.n939 VPWR.n327 0.369731
R4468 VPWR.n941 VPWR.n940 0.369731
R4469 VPWR.n945 VPWR.n325 0.369731
R4470 VPWR.n947 VPWR.n946 0.369731
R4471 VPWR.n972 VPWR.n314 0.369731
R4472 VPWR.n974 VPWR.n973 0.369731
R4473 VPWR.n978 VPWR.n312 0.369731
R4474 VPWR.n733 VPWR.n439 0.369731
R4475 VPWR.n761 VPWR.n759 0.369731
R4476 VPWR.n710 VPWR.n695 0.369731
R4477 VPWR.n728 VPWR.n727 0.369731
R4478 VPWR.n521 VPWR.n520 0.369731
R4479 VPWR.n678 VPWR.n677 0.369731
R4480 VPWR.n26 VPWR.n4 0.318338
R4481 VPWR.n102 VPWR.n80 0.318338
R4482 VPWR.n43 VPWR.n40 0.305262
R4483 VPWR.n1129 VPWR.n1128 0.305262
R4484 VPWR.n1122 VPWR.n50 0.305262
R4485 VPWR.n1118 VPWR.n1117 0.305262
R4486 VPWR.n786 VPWR.n778 0.305262
R4487 VPWR.n839 VPWR.n800 0.305262
R4488 VPWR.n824 VPWR.n815 0.305262
R4489 VPWR.n473 VPWR.n472 0.305262
R4490 VPWR.n547 VPWR.n460 0.305262
R4491 VPWR.n163 VPWR.n162 0.305262
R4492 VPWR.n170 VPWR.n169 0.305262
R4493 VPWR.n162 VPWR.n161 0.254468
R4494 VPWR.n904 VPWR 0.238178
R4495 VPWR.n427 VPWR 0.238178
R4496 VPWR.n397 VPWR.n396 0.227049
R4497 VPWR.n384 VPWR.n366 0.227049
R4498 VPWR.n984 VPWR.n983 0.227049
R4499 VPWR.n1004 VPWR.n1003 0.227049
R4500 VPWR.n555 VPWR.n554 0.227049
R4501 VPWR.n644 VPWR.n643 0.227049
R4502 VPWR.n102 VPWR.n26 0.2167
R4503 VPWR.n1189 VPWR.n8 0.21207
R4504 VPWR.n1177 VPWR.n15 0.21207
R4505 VPWR.n777 VPWR.n776 0.203675
R4506 VPWR.n861 VPWR.n860 0.203675
R4507 VPWR.n904 VPWR.n890 0.19052
R4508 VPWR.n427 VPWR.n415 0.19052
R4509 VPWR.n1086 VPWR 0.17983
R4510 VPWR VPWR.n1054 0.17983
R4511 VPWR.n822 VPWR 0.17983
R4512 VPWR VPWR.n612 0.17983
R4513 VPWR VPWR.n240 0.17983
R4514 VPWR VPWR.n1055 0.179485
R4515 VPWR.n138 VPWR 0.179485
R4516 VPWR VPWR.n354 0.172576
R4517 VPWR VPWR.n903 0.172576
R4518 VPWR VPWR.n426 0.172576
R4519 VPWR VPWR.n470 0.172576
R4520 VPWR.n156 VPWR 0.172576
R4521 VPWR.n536 VPWR.n535 0.163904
R4522 VPWR.n527 VPWR.n526 0.163904
R4523 VPWR.n306 VPWR.n290 0.1603
R4524 VPWR.n995 VPWR.n306 0.1603
R4525 VPWR.n995 VPWR.n307 0.1603
R4526 VPWR.n572 VPWR.n307 0.1603
R4527 VPWR.n1161 VPWR.n1160 0.1603
R4528 VPWR.n1160 VPWR.n29 0.1603
R4529 VPWR.n739 VPWR.n29 0.1603
R4530 VPWR.n739 VPWR.n684 0.1603
R4531 VPWR.n411 VPWR.n4 0.1603
R4532 VPWR.n915 VPWR.n411 0.1603
R4533 VPWR.n915 VPWR.n888 0.1603
R4534 VPWR.n888 VPWR.n413 0.1603
R4535 VPWR.n1074 VPWR.n80 0.1603
R4536 VPWR.n1074 VPWR.n1065 0.1603
R4537 VPWR.n1065 VPWR.n82 0.1603
R4538 VPWR.n599 VPWR.n82 0.1603
R4539 VPWR.n1055 VPWR 0.14207
R4540 VPWR.n1086 VPWR 0.141725
R4541 VPWR.n1054 VPWR 0.141725
R4542 VPWR.n822 VPWR 0.141725
R4543 VPWR.n612 VPWR 0.141725
R4544 VPWR.n240 VPWR 0.141725
R4545 VPWR VPWR.n138 0.140768
R4546 VPWR.n355 VPWR 0.120408
R4547 VPWR.n356 VPWR 0.120408
R4548 VPWR.n398 VPWR.n363 0.120292
R4549 VPWR.n392 VPWR.n363 0.120292
R4550 VPWR.n392 VPWR.n391 0.120292
R4551 VPWR.n391 VPWR.n390 0.120292
R4552 VPWR.n390 VPWR.n365 0.120292
R4553 VPWR.n386 VPWR.n365 0.120292
R4554 VPWR.n386 VPWR.n385 0.120292
R4555 VPWR.n382 VPWR.n381 0.120292
R4556 VPWR.n381 VPWR.n368 0.120292
R4557 VPWR.n376 VPWR.n368 0.120292
R4558 VPWR.n376 VPWR.n375 0.120292
R4559 VPWR.n375 VPWR.n371 0.120292
R4560 VPWR.n1144 VPWR.n37 0.120292
R4561 VPWR.n1139 VPWR.n37 0.120292
R4562 VPWR.n1139 VPWR.n1138 0.120292
R4563 VPWR.n1134 VPWR.n1133 0.120292
R4564 VPWR.n1133 VPWR.n41 0.120292
R4565 VPWR.n1127 VPWR.n41 0.120292
R4566 VPWR.n1121 VPWR.n1120 0.120292
R4567 VPWR.n1120 VPWR.n51 0.120292
R4568 VPWR.n1112 VPWR.n58 0.120292
R4569 VPWR.n60 VPWR.n58 0.120292
R4570 VPWR.n1107 VPWR.n60 0.120292
R4571 VPWR.n1105 VPWR.n63 0.120292
R4572 VPWR.n67 VPWR.n64 0.120292
R4573 VPWR.n68 VPWR.n67 0.120292
R4574 VPWR.n1099 VPWR.n68 0.120292
R4575 VPWR.n1098 VPWR.n1097 0.120292
R4576 VPWR.n1092 VPWR.n1091 0.120292
R4577 VPWR.n1091 VPWR.n1090 0.120292
R4578 VPWR.n1090 VPWR.n1078 0.120292
R4579 VPWR.n926 VPWR.n925 0.120292
R4580 VPWR.n926 VPWR.n330 0.120292
R4581 VPWR.n931 VPWR.n330 0.120292
R4582 VPWR.n932 VPWR.n931 0.120292
R4583 VPWR.n933 VPWR.n932 0.120292
R4584 VPWR.n933 VPWR.n328 0.120292
R4585 VPWR.n937 VPWR.n328 0.120292
R4586 VPWR.n938 VPWR.n937 0.120292
R4587 VPWR.n943 VPWR.n326 0.120292
R4588 VPWR.n944 VPWR.n943 0.120292
R4589 VPWR.n964 VPWR.n317 0.120292
R4590 VPWR.n965 VPWR.n964 0.120292
R4591 VPWR.n966 VPWR.n965 0.120292
R4592 VPWR.n966 VPWR.n315 0.120292
R4593 VPWR.n970 VPWR.n315 0.120292
R4594 VPWR.n971 VPWR.n970 0.120292
R4595 VPWR.n976 VPWR.n313 0.120292
R4596 VPWR.n977 VPWR.n976 0.120292
R4597 VPWR.n986 VPWR.n309 0.120292
R4598 VPWR.n1005 VPWR.n96 0.120292
R4599 VPWR.n1011 VPWR.n1010 0.120292
R4600 VPWR.n1012 VPWR.n1011 0.120292
R4601 VPWR.n1017 VPWR.n1016 0.120292
R4602 VPWR.n1017 VPWR.n90 0.120292
R4603 VPWR.n1021 VPWR.n90 0.120292
R4604 VPWR.n1022 VPWR.n1021 0.120292
R4605 VPWR.n1028 VPWR.n87 0.120292
R4606 VPWR.n1029 VPWR.n1028 0.120292
R4607 VPWR.n712 VPWR.n711 0.120292
R4608 VPWR.n712 VPWR.n694 0.120292
R4609 VPWR.n717 VPWR.n694 0.120292
R4610 VPWR.n718 VPWR.n717 0.120292
R4611 VPWR.n718 VPWR.n692 0.120292
R4612 VPWR.n722 VPWR.n692 0.120292
R4613 VPWR.n723 VPWR.n722 0.120292
R4614 VPWR.n724 VPWR.n723 0.120292
R4615 VPWR.n724 VPWR.n690 0.120292
R4616 VPWR.n729 VPWR.n690 0.120292
R4617 VPWR.n749 VPWR.n438 0.120292
R4618 VPWR.n750 VPWR.n749 0.120292
R4619 VPWR.n750 VPWR.n436 0.120292
R4620 VPWR.n754 VPWR.n436 0.120292
R4621 VPWR.n755 VPWR.n754 0.120292
R4622 VPWR.n756 VPWR.n755 0.120292
R4623 VPWR.n756 VPWR.n434 0.120292
R4624 VPWR.n762 VPWR.n434 0.120292
R4625 VPWR.n864 VPWR.n863 0.120292
R4626 VPWR.n863 VPWR.n785 0.120292
R4627 VPWR.n856 VPWR.n855 0.120292
R4628 VPWR.n851 VPWR.n850 0.120292
R4629 VPWR.n850 VPWR.n849 0.120292
R4630 VPWR.n849 VPWR.n794 0.120292
R4631 VPWR.n844 VPWR.n843 0.120292
R4632 VPWR.n843 VPWR.n842 0.120292
R4633 VPWR.n827 VPWR.n826 0.120292
R4634 VPWR.n826 VPWR.n825 0.120292
R4635 VPWR.n477 VPWR.n461 0.120292
R4636 VPWR.n537 VPWR.n486 0.120292
R4637 VPWR.n531 VPWR.n486 0.120292
R4638 VPWR.n531 VPWR.n530 0.120292
R4639 VPWR.n530 VPWR.n529 0.120292
R4640 VPWR.n529 VPWR.n492 0.120292
R4641 VPWR.n522 VPWR.n494 0.120292
R4642 VPWR.n517 VPWR.n494 0.120292
R4643 VPWR.n517 VPWR.n516 0.120292
R4644 VPWR.n516 VPWR.n496 0.120292
R4645 VPWR.n511 VPWR.n496 0.120292
R4646 VPWR.n511 VPWR.n510 0.120292
R4647 VPWR.n680 VPWR.n449 0.120292
R4648 VPWR.n670 VPWR.n669 0.120292
R4649 VPWR.n668 VPWR.n454 0.120292
R4650 VPWR.n663 VPWR.n454 0.120292
R4651 VPWR.n663 VPWR.n662 0.120292
R4652 VPWR.n658 VPWR.n657 0.120292
R4653 VPWR.n649 VPWR.n648 0.120292
R4654 VPWR.n648 VPWR.n647 0.120292
R4655 VPWR.n647 VPWR.n576 0.120292
R4656 VPWR.n642 VPWR.n576 0.120292
R4657 VPWR.n641 VPWR.n640 0.120292
R4658 VPWR.n640 VPWR.n579 0.120292
R4659 VPWR.n636 VPWR.n635 0.120292
R4660 VPWR.n631 VPWR.n583 0.120292
R4661 VPWR.n631 VPWR.n630 0.120292
R4662 VPWR.n630 VPWR.n629 0.120292
R4663 VPWR.n618 VPWR.n601 0.120292
R4664 VPWR.n614 VPWR.n601 0.120292
R4665 VPWR.n614 VPWR.n613 0.120292
R4666 VPWR.n165 VPWR.n164 0.120292
R4667 VPWR.n165 VPWR.n150 0.120292
R4668 VPWR.n171 VPWR.n150 0.120292
R4669 VPWR.n1188 VPWR.n1187 0.120292
R4670 VPWR.n1187 VPWR.n9 0.120292
R4671 VPWR.n1182 VPWR.n9 0.120292
R4672 VPWR.n1181 VPWR.n13 0.120292
R4673 VPWR.n1176 VPWR.n13 0.120292
R4674 VPWR.n1176 VPWR.n1175 0.120292
R4675 VPWR.n1175 VPWR.n16 0.120292
R4676 VPWR.n1170 VPWR.n16 0.120292
R4677 VPWR.n1169 VPWR.n1168 0.120292
R4678 VPWR.n115 VPWR.n112 0.120292
R4679 VPWR.n146 VPWR.n145 0.120292
R4680 VPWR.n200 VPWR.n197 0.120292
R4681 VPWR.n273 VPWR.n205 0.120292
R4682 VPWR.n266 VPWR.n205 0.120292
R4683 VPWR.n259 VPWR.n258 0.120292
R4684 VPWR.n246 VPWR.n229 0.120292
R4685 VPWR.n242 VPWR.n229 0.120292
R4686 VPWR.n242 VPWR.n241 0.120292
R4687 VPWR.n651 VPWR.n556 0.113774
R4688 VPWR.n354 VPWR 0.105238
R4689 VPWR.n903 VPWR 0.105238
R4690 VPWR.n426 VPWR 0.105238
R4691 VPWR.n470 VPWR 0.105238
R4692 VPWR.n156 VPWR 0.105238
R4693 VPWR.n290 VPWR.n102 0.102137
R4694 VPWR.n1161 VPWR.n26 0.102137
R4695 VPWR.n776 VPWR.n775 0.102087
R4696 VPWR.n860 VPWR.n787 0.102087
R4697 VPWR.n168 VPWR.n167 0.102087
R4698 VPWR VPWR.n326 0.0981562
R4699 VPWR VPWR.n313 0.0981562
R4700 VPWR.n980 VPWR 0.0981562
R4701 VPWR.n1010 VPWR 0.0981562
R4702 VPWR.n730 VPWR 0.0981562
R4703 VPWR.n763 VPWR 0.0981562
R4704 VPWR.n764 VPWR 0.0981562
R4705 VPWR VPWR.n461 0.0981562
R4706 VPWR.n674 VPWR 0.0981562
R4707 VPWR VPWR.n673 0.0981562
R4708 VPWR.n670 VPWR 0.0981562
R4709 VPWR.n583 VPWR 0.0981562
R4710 VPWR.n1165 VPWR 0.0981562
R4711 VPWR.n185 VPWR 0.0981562
R4712 VPWR VPWR.n278 0.0981562
R4713 VPWR VPWR.n273 0.0981562
R4714 VPWR VPWR.n264 0.0981562
R4715 VPWR VPWR.n259 0.0981562
R4716 VPWR VPWR.n1105 0.0968542
R4717 VPWR.n175 VPWR.n174 0.0950946
R4718 VPWR.n1193 VPWR.n2 0.0950946
R4719 VPWR.n1163 VPWR.n24 0.0950946
R4720 VPWR.n132 VPWR.n131 0.0950946
R4721 VPWR.n288 VPWR.n287 0.0950946
R4722 VPWR.n195 VPWR.n194 0.0950946
R4723 VPWR.n1158 VPWR.n1157 0.0950946
R4724 VPWR.n1150 VPWR.n1149 0.0950946
R4725 VPWR.n409 VPWR.n408 0.0950946
R4726 VPWR.n401 VPWR.n400 0.0950946
R4727 VPWR.n1072 VPWR.n1071 0.0950946
R4728 VPWR.n1076 VPWR.n78 0.0950946
R4729 VPWR.n304 VPWR.n303 0.0950946
R4730 VPWR.n296 VPWR.n294 0.0950946
R4731 VPWR.n951 VPWR.n950 0.0950946
R4732 VPWR.n957 VPWR.n956 0.0950946
R4733 VPWR.n913 VPWR.n912 0.0950946
R4734 VPWR.n918 VPWR.n917 0.0950946
R4735 VPWR.n1063 VPWR.n1062 0.0950946
R4736 VPWR.n1045 VPWR.n1044 0.0950946
R4737 VPWR.n993 VPWR.n992 0.0950946
R4738 VPWR.n998 VPWR.n997 0.0950946
R4739 VPWR.n570 VPWR.n569 0.0950946
R4740 VPWR.n574 VPWR.n559 0.0950946
R4741 VPWR.n873 VPWR.n768 0.0950946
R4742 VPWR.n783 VPWR.n780 0.0950946
R4743 VPWR.n886 VPWR.n885 0.0950946
R4744 VPWR.n703 VPWR.n702 0.0950946
R4745 VPWR.n806 VPWR.n805 0.0950946
R4746 VPWR.n832 VPWR.n804 0.0950946
R4747 VPWR.n737 VPWR.n736 0.0950946
R4748 VPWR.n742 VPWR.n741 0.0950946
R4749 VPWR.n508 VPWR.n507 0.0950946
R4750 VPWR.n682 VPWR.n447 0.0950946
R4751 VPWR.n597 VPWR.n596 0.0950946
R4752 VPWR.n620 VPWR.n594 0.0950946
R4753 VPWR.n544 VPWR.n479 0.0950946
R4754 VPWR.n539 VPWR.n482 0.0950946
R4755 VPWR.n224 VPWR.n223 0.0950946
R4756 VPWR.n248 VPWR.n221 0.0950946
R4757 VPWR VPWR.n355 0.0930646
R4758 VPWR.n572 VPWR 0.08745
R4759 VPWR.n684 VPWR 0.08745
R4760 VPWR.n413 VPWR 0.08745
R4761 VPWR.n599 VPWR 0.08745
R4762 VPWR.n1151 VPWR.n1145 0.0838333
R4763 VPWR.n1077 VPWR.n77 0.0838333
R4764 VPWR.n919 VPWR.n334 0.0838333
R4765 VPWR.n958 VPWR.n320 0.0838333
R4766 VPWR.n991 VPWR.n987 0.0838333
R4767 VPWR.n999 VPWR.n99 0.0838333
R4768 VPWR.n1046 VPWR.n1039 0.0838333
R4769 VPWR.n704 VPWR.n697 0.0838333
R4770 VPWR.n743 VPWR.n441 0.0838333
R4771 VPWR.n831 VPWR.n809 0.0838333
R4772 VPWR.n509 VPWR.n498 0.0838333
R4773 VPWR.n681 VPWR.n448 0.0838333
R4774 VPWR.n575 VPWR.n558 0.0838333
R4775 VPWR.n619 VPWR.n600 0.0838333
R4776 VPWR.n196 VPWR.n190 0.0838333
R4777 VPWR.n247 VPWR.n228 0.0838333
R4778 VPWR.n332 VPWR 0.082648
R4779 VPWR.n949 VPWR 0.0747188
R4780 VPWR.n1061 VPWR 0.0747188
R4781 VPWR.n735 VPWR 0.0747188
R4782 VPWR.n568 VPWR 0.0747188
R4783 VPWR.n124 VPWR 0.0747188
R4784 VPWR.n356 VPWR.n339 0.0735334
R4785 VPWR.n334 VPWR.n332 0.0735334
R4786 VPWR.n1197 VPWR.n1 0.0680676
R4787 VPWR.n1197 VPWR.n1196 0.0680676
R4788 VPWR.n128 VPWR.n127 0.0680676
R4789 VPWR.n130 VPWR.n128 0.0680676
R4790 VPWR.n191 VPWR.n106 0.0680676
R4791 VPWR.n193 VPWR.n191 0.0680676
R4792 VPWR.n1146 VPWR.n32 0.0680676
R4793 VPWR.n1148 VPWR.n1146 0.0680676
R4794 VPWR.n360 VPWR.n340 0.0680676
R4795 VPWR.n362 VPWR.n360 0.0680676
R4796 VPWR.n1069 VPWR.n1068 0.0680676
R4797 VPWR.n1068 VPWR.n1067 0.0680676
R4798 VPWR.n301 VPWR.n300 0.0680676
R4799 VPWR.n300 VPWR.n298 0.0680676
R4800 VPWR.n323 VPWR.n322 0.0680676
R4801 VPWR.n322 VPWR.n321 0.0680676
R4802 VPWR.n892 VPWR.n891 0.0680676
R4803 VPWR.n891 VPWR.n335 0.0680676
R4804 VPWR.n1041 VPWR.n85 0.0680676
R4805 VPWR.n1043 VPWR.n1041 0.0680676
R4806 VPWR.n989 VPWR.n988 0.0680676
R4807 VPWR.n988 VPWR.n100 0.0680676
R4808 VPWR.n565 VPWR.n562 0.0680676
R4809 VPWR.n565 VPWR.n564 0.0680676
R4810 VPWR.n870 VPWR.n869 0.0680676
R4811 VPWR.n869 VPWR.n770 0.0680676
R4812 VPWR.n699 VPWR.n416 0.0680676
R4813 VPWR.n701 VPWR.n699 0.0680676
R4814 VPWR.n836 VPWR.n803 0.0680676
R4815 VPWR.n836 VPWR.n835 0.0680676
R4816 VPWR.n688 VPWR.n687 0.0680676
R4817 VPWR.n687 VPWR.n442 0.0680676
R4818 VPWR.n506 VPWR.n504 0.0680676
R4819 VPWR.n504 VPWR.n499 0.0680676
R4820 VPWR.n624 VPWR.n593 0.0680676
R4821 VPWR.n624 VPWR.n623 0.0680676
R4822 VPWR.n483 VPWR.n480 0.0680676
R4823 VPWR.n483 VPWR.n481 0.0680676
R4824 VPWR.n252 VPWR.n220 0.0680676
R4825 VPWR.n252 VPWR.n251 0.0680676
R4826 VPWR.n403 VPWR 0.0603958
R4827 VPWR.n382 VPWR 0.0603958
R4828 VPWR.n1155 VPWR.n33 0.0603958
R4829 VPWR.n1152 VPWR.n33 0.0603958
R4830 VPWR.n1135 VPWR 0.0603958
R4831 VPWR VPWR.n1134 0.0603958
R4832 VPWR VPWR.n1126 0.0603958
R4833 VPWR VPWR.n1125 0.0603958
R4834 VPWR.n1121 VPWR 0.0603958
R4835 VPWR.n299 VPWR.n54 0.0603958
R4836 VPWR VPWR.n1112 0.0603958
R4837 VPWR.n1107 VPWR 0.0603958
R4838 VPWR VPWR.n1106 0.0603958
R4839 VPWR.n64 VPWR 0.0603958
R4840 VPWR.n1099 VPWR 0.0603958
R4841 VPWR VPWR.n1098 0.0603958
R4842 VPWR VPWR.n73 0.0603958
R4843 VPWR VPWR.n1078 0.0603958
R4844 VPWR.n920 VPWR 0.0603958
R4845 VPWR.n925 VPWR 0.0603958
R4846 VPWR.n948 VPWR.n319 0.0603958
R4847 VPWR.n959 VPWR.n319 0.0603958
R4848 VPWR.n981 VPWR 0.0603958
R4849 VPWR VPWR.n309 0.0603958
R4850 VPWR.n990 VPWR.n98 0.0603958
R4851 VPWR.n1000 VPWR.n98 0.0603958
R4852 VPWR.n1006 VPWR 0.0603958
R4853 VPWR.n1016 VPWR 0.0603958
R4854 VPWR VPWR.n87 0.0603958
R4855 VPWR.n1040 VPWR.n1031 0.0603958
R4856 VPWR VPWR.n698 0.0603958
R4857 VPWR.n707 VPWR 0.0603958
R4858 VPWR.n711 VPWR 0.0603958
R4859 VPWR.n734 VPWR.n440 0.0603958
R4860 VPWR.n744 VPWR.n440 0.0603958
R4861 VPWR.n766 VPWR 0.0603958
R4862 VPWR.n875 VPWR 0.0603958
R4863 VPWR.n868 VPWR.n772 0.0603958
R4864 VPWR.n868 VPWR 0.0603958
R4865 VPWR VPWR.n864 0.0603958
R4866 VPWR VPWR.n856 0.0603958
R4867 VPWR.n855 VPWR 0.0603958
R4868 VPWR.n851 VPWR 0.0603958
R4869 VPWR.n844 VPWR 0.0603958
R4870 VPWR.n838 VPWR.n837 0.0603958
R4871 VPWR.n837 VPWR.n802 0.0603958
R4872 VPWR.n827 VPWR 0.0603958
R4873 VPWR.n471 VPWR 0.0603958
R4874 VPWR VPWR.n477 0.0603958
R4875 VPWR.n546 VPWR 0.0603958
R4876 VPWR.n484 VPWR 0.0603958
R4877 VPWR.n523 VPWR 0.0603958
R4878 VPWR VPWR.n522 0.0603958
R4879 VPWR.n503 VPWR.n501 0.0603958
R4880 VPWR.n503 VPWR.n502 0.0603958
R4881 VPWR.n669 VPWR 0.0603958
R4882 VPWR VPWR.n668 0.0603958
R4883 VPWR VPWR.n661 0.0603958
R4884 VPWR.n658 VPWR 0.0603958
R4885 VPWR VPWR.n656 0.0603958
R4886 VPWR.n567 VPWR.n566 0.0603958
R4887 VPWR.n566 VPWR.n563 0.0603958
R4888 VPWR VPWR.n641 0.0603958
R4889 VPWR VPWR.n579 0.0603958
R4890 VPWR.n636 VPWR 0.0603958
R4891 VPWR.n625 VPWR.n592 0.0603958
R4892 VPWR.n613 VPWR 0.0603958
R4893 VPWR.n164 VPWR 0.0603958
R4894 VPWR VPWR.n0 0.0603958
R4895 VPWR.n1188 VPWR 0.0603958
R4896 VPWR VPWR.n1181 0.0603958
R4897 VPWR VPWR.n1169 0.0603958
R4898 VPWR.n126 VPWR.n125 0.0603958
R4899 VPWR.n134 VPWR.n126 0.0603958
R4900 VPWR.n139 VPWR 0.0603958
R4901 VPWR VPWR.n115 0.0603958
R4902 VPWR.n112 VPWR 0.0603958
R4903 VPWR VPWR.n111 0.0603958
R4904 VPWR.n145 VPWR 0.0603958
R4905 VPWR.n147 VPWR 0.0603958
R4906 VPWR.n183 VPWR 0.0603958
R4907 VPWR.n184 VPWR 0.0603958
R4908 VPWR VPWR.n189 0.0603958
R4909 VPWR VPWR.n200 0.0603958
R4910 VPWR.n279 VPWR 0.0603958
R4911 VPWR.n278 VPWR 0.0603958
R4912 VPWR.n274 VPWR 0.0603958
R4913 VPWR.n266 VPWR 0.0603958
R4914 VPWR VPWR.n265 0.0603958
R4915 VPWR.n264 VPWR 0.0603958
R4916 VPWR.n260 VPWR 0.0603958
R4917 VPWR.n258 VPWR 0.0603958
R4918 VPWR.n214 VPWR 0.0603958
R4919 VPWR.n253 VPWR.n219 0.0603958
R4920 VPWR.n241 VPWR 0.0603958
R4921 VPWR.n1195 VPWR.n3 0.0574697
R4922 VPWR.n129 VPWR.n25 0.0574697
R4923 VPWR.n192 VPWR.n104 0.0574697
R4924 VPWR.n1147 VPWR.n30 0.0574697
R4925 VPWR.n361 VPWR.n338 0.0574697
R4926 VPWR.n1066 VPWR.n79 0.0574697
R4927 VPWR.n297 VPWR.n292 0.0574697
R4928 VPWR.n954 VPWR.n953 0.0574697
R4929 VPWR.n889 VPWR.n336 0.0574697
R4930 VPWR.n1042 VPWR.n83 0.0574697
R4931 VPWR.n308 VPWR.n101 0.0574697
R4932 VPWR.n561 VPWR.n560 0.0574697
R4933 VPWR.n872 VPWR.n871 0.0574697
R4934 VPWR.n782 VPWR.n781 0.0574697
R4935 VPWR.n700 VPWR.n414 0.0574697
R4936 VPWR.n834 VPWR.n808 0.0574697
R4937 VPWR.n685 VPWR.n443 0.0574697
R4938 VPWR.n505 VPWR.n445 0.0574697
R4939 VPWR.n683 VPWR.n446 0.0574697
R4940 VPWR.n622 VPWR.n595 0.0574697
R4941 VPWR.n542 VPWR.n541 0.0574697
R4942 VPWR.n226 VPWR.n225 0.0574697
R4943 VPWR.n250 VPWR.n249 0.0574697
R4944 VPWR.n534 VPWR.n533 0.0549681
R4945 VPWR.n399 VPWR 0.047375
R4946 VPWR VPWR.n57 0.047375
R4947 VPWR.n784 VPWR 0.047375
R4948 VPWR.n538 VPWR 0.047375
R4949 VPWR.n1192 VPWR 0.047375
R4950 VPWR VPWR.n122 0.047375
R4951 VPWR VPWR.n105 0.047375
R4952 VPWR.n175 VPWR.n1 0.0410405
R4953 VPWR.n1196 VPWR.n2 0.0410405
R4954 VPWR.n127 VPWR.n24 0.0410405
R4955 VPWR.n132 VPWR.n130 0.0410405
R4956 VPWR.n287 VPWR.n106 0.0410405
R4957 VPWR.n194 VPWR.n193 0.0410405
R4958 VPWR.n1157 VPWR.n32 0.0410405
R4959 VPWR.n1150 VPWR.n1148 0.0410405
R4960 VPWR.n408 VPWR.n340 0.0410405
R4961 VPWR.n401 VPWR.n362 0.0410405
R4962 VPWR.n1071 VPWR.n1069 0.0410405
R4963 VPWR.n1067 VPWR.n78 0.0410405
R4964 VPWR.n303 VPWR.n301 0.0410405
R4965 VPWR.n298 VPWR.n296 0.0410405
R4966 VPWR.n950 VPWR.n323 0.0410405
R4967 VPWR.n957 VPWR.n321 0.0410405
R4968 VPWR.n912 VPWR.n892 0.0410405
R4969 VPWR.n918 VPWR.n335 0.0410405
R4970 VPWR.n1062 VPWR.n85 0.0410405
R4971 VPWR.n1044 VPWR.n1043 0.0410405
R4972 VPWR.n992 VPWR.n989 0.0410405
R4973 VPWR.n998 VPWR.n100 0.0410405
R4974 VPWR.n569 VPWR.n562 0.0410405
R4975 VPWR.n564 VPWR.n559 0.0410405
R4976 VPWR.n870 VPWR.n768 0.0410405
R4977 VPWR.n780 VPWR.n770 0.0410405
R4978 VPWR.n885 VPWR.n416 0.0410405
R4979 VPWR.n702 VPWR.n701 0.0410405
R4980 VPWR.n805 VPWR.n803 0.0410405
R4981 VPWR.n835 VPWR.n804 0.0410405
R4982 VPWR.n736 VPWR.n688 0.0410405
R4983 VPWR.n742 VPWR.n442 0.0410405
R4984 VPWR.n507 VPWR.n506 0.0410405
R4985 VPWR.n499 VPWR.n447 0.0410405
R4986 VPWR.n596 VPWR.n593 0.0410405
R4987 VPWR.n623 VPWR.n594 0.0410405
R4988 VPWR.n480 VPWR.n479 0.0410405
R4989 VPWR.n482 VPWR.n481 0.0410405
R4990 VPWR.n223 VPWR.n220 0.0410405
R4991 VPWR.n251 VPWR.n221 0.0410405
R4992 VPWR.n1040 VPWR 0.0382604
R4993 VPWR VPWR.n625 0.0382604
R4994 VPWR VPWR.n253 0.0382604
R4995 VPWR.n407 VPWR 0.0369583
R4996 VPWR.n1156 VPWR 0.0369583
R4997 VPWR.n302 VPWR 0.0369583
R4998 VPWR.n299 VPWR 0.0369583
R4999 VPWR.n295 VPWR 0.0369583
R5000 VPWR.n1070 VPWR 0.0369583
R5001 VPWR.n911 VPWR 0.0369583
R5002 VPWR.n884 VPWR 0.0369583
R5003 VPWR.n771 VPWR 0.0369583
R5004 VPWR.n779 VPWR 0.0369583
R5005 VPWR.n801 VPWR 0.0369583
R5006 VPWR.n478 VPWR 0.0369583
R5007 VPWR.n591 VPWR 0.0369583
R5008 VPWR.n176 VPWR 0.0369583
R5009 VPWR VPWR.n5 0.0369583
R5010 VPWR.n133 VPWR 0.0369583
R5011 VPWR.n286 VPWR 0.0369583
R5012 VPWR VPWR.n218 0.0369583
R5013 VPWR VPWR.n706 0.0330521
R5014 VPWR.n657 VPWR 0.0330521
R5015 VPWR VPWR.n146 0.0330521
R5016 VPWR.n406 VPWR 0.03175
R5017 VPWR.n1135 VPWR 0.03175
R5018 VPWR.n1125 VPWR 0.03175
R5019 VPWR.n1113 VPWR 0.03175
R5020 VPWR.n910 VPWR 0.03175
R5021 VPWR VPWR.n980 0.03175
R5022 VPWR.n981 VPWR 0.03175
R5023 VPWR.n883 VPWR 0.03175
R5024 VPWR VPWR.n764 0.03175
R5025 VPWR VPWR.n766 0.03175
R5026 VPWR.n865 VPWR 0.03175
R5027 VPWR VPWR.n459 0.03175
R5028 VPWR.n661 VPWR 0.03175
R5029 VPWR.n177 VPWR 0.03175
R5030 VPWR.n1191 VPWR 0.03175
R5031 VPWR.n147 VPWR 0.03175
R5032 VPWR.n571 VPWR.n561 0.0292489
R5033 VPWR.n573 VPWR.n560 0.0292489
R5034 VPWR.n994 VPWR.n308 0.0292489
R5035 VPWR.n996 VPWR.n101 0.0292489
R5036 VPWR.n305 VPWR.n292 0.0292489
R5037 VPWR.n297 VPWR.n291 0.0292489
R5038 VPWR.n289 VPWR.n104 0.0292489
R5039 VPWR.n192 VPWR.n103 0.0292489
R5040 VPWR.n781 VPWR.n769 0.0292489
R5041 VPWR.n871 VPWR.n769 0.0292489
R5042 VPWR.n738 VPWR.n685 0.0292489
R5043 VPWR.n740 VPWR.n443 0.0292489
R5044 VPWR.n953 VPWR.n952 0.0292489
R5045 VPWR.n955 VPWR.n954 0.0292489
R5046 VPWR.n1159 VPWR.n30 0.0292489
R5047 VPWR.n1147 VPWR.n28 0.0292489
R5048 VPWR.n1162 VPWR.n25 0.0292489
R5049 VPWR.n129 VPWR.n27 0.0292489
R5050 VPWR.n446 VPWR.n444 0.0292489
R5051 VPWR.n505 VPWR.n444 0.0292489
R5052 VPWR.n543 VPWR.n542 0.0292489
R5053 VPWR.n541 VPWR.n540 0.0292489
R5054 VPWR.n887 VPWR.n414 0.0292489
R5055 VPWR.n700 VPWR.n412 0.0292489
R5056 VPWR.n914 VPWR.n889 0.0292489
R5057 VPWR.n916 VPWR.n336 0.0292489
R5058 VPWR.n410 VPWR.n338 0.0292489
R5059 VPWR.n361 VPWR.n337 0.0292489
R5060 VPWR.n173 VPWR.n3 0.0292489
R5061 VPWR.n1195 VPWR.n1194 0.0292489
R5062 VPWR.n598 VPWR.n595 0.0292489
R5063 VPWR.n622 VPWR.n621 0.0292489
R5064 VPWR.n808 VPWR.n807 0.0292489
R5065 VPWR.n834 VPWR.n833 0.0292489
R5066 VPWR.n1064 VPWR.n83 0.0292489
R5067 VPWR.n1042 VPWR.n81 0.0292489
R5068 VPWR.n1073 VPWR.n1066 0.0292489
R5069 VPWR.n1075 VPWR.n79 0.0292489
R5070 VPWR.n250 VPWR.n227 0.0292489
R5071 VPWR.n227 VPWR.n226 0.0292489
R5072 VPWR.n407 VPWR.n406 0.0239375
R5073 VPWR.n403 VPWR.n402 0.0239375
R5074 VPWR.n1156 VPWR.n1155 0.0239375
R5075 VPWR.n1152 VPWR.n1151 0.0239375
R5076 VPWR.n302 VPWR.n53 0.0239375
R5077 VPWR VPWR.n53 0.0239375
R5078 VPWR.n1106 VPWR 0.0239375
R5079 VPWR.n1070 VPWR.n72 0.0239375
R5080 VPWR.n911 VPWR.n910 0.0239375
R5081 VPWR.n920 VPWR.n919 0.0239375
R5082 VPWR.n949 VPWR.n948 0.0239375
R5083 VPWR.n959 VPWR.n958 0.0239375
R5084 VPWR.n991 VPWR.n990 0.0239375
R5085 VPWR.n1000 VPWR.n999 0.0239375
R5086 VPWR.n1061 VPWR.n1060 0.0239375
R5087 VPWR.n1039 VPWR.n1031 0.0239375
R5088 VPWR.n884 VPWR.n883 0.0239375
R5089 VPWR.n698 VPWR.n697 0.0239375
R5090 VPWR.n735 VPWR.n734 0.0239375
R5091 VPWR.n744 VPWR.n743 0.0239375
R5092 VPWR.n772 VPWR.n771 0.0239375
R5093 VPWR.n838 VPWR.n801 0.0239375
R5094 VPWR.n809 VPWR.n802 0.0239375
R5095 VPWR.n478 VPWR.n459 0.0239375
R5096 VPWR.n485 VPWR.n484 0.0239375
R5097 VPWR.n501 VPWR.n498 0.0239375
R5098 VPWR.n502 VPWR.n448 0.0239375
R5099 VPWR.n568 VPWR.n567 0.0239375
R5100 VPWR.n563 VPWR.n558 0.0239375
R5101 VPWR.n626 VPWR.n591 0.0239375
R5102 VPWR.n600 VPWR.n592 0.0239375
R5103 VPWR.n177 VPWR.n176 0.0239375
R5104 VPWR.n125 VPWR.n124 0.0239375
R5105 VPWR.n134 VPWR.n133 0.0239375
R5106 VPWR.n286 VPWR.n285 0.0239375
R5107 VPWR.n254 VPWR.n218 0.0239375
R5108 VPWR.n228 VPWR.n219 0.0239375
R5109 VPWR.n385 VPWR 0.0226354
R5110 VPWR.n1138 VPWR 0.0226354
R5111 VPWR.n1127 VPWR 0.0226354
R5112 VPWR.n1126 VPWR 0.0226354
R5113 VPWR VPWR.n54 0.0226354
R5114 VPWR VPWR.n63 0.0226354
R5115 VPWR VPWR.n72 0.0226354
R5116 VPWR.n938 VPWR 0.0226354
R5117 VPWR.n971 VPWR 0.0226354
R5118 VPWR.n977 VPWR 0.0226354
R5119 VPWR VPWR.n1005 0.0226354
R5120 VPWR.n1006 VPWR 0.0226354
R5121 VPWR.n1012 VPWR 0.0226354
R5122 VPWR.n1022 VPWR 0.0226354
R5123 VPWR.n1060 VPWR 0.0226354
R5124 VPWR.n1056 VPWR 0.0226354
R5125 VPWR.n707 VPWR 0.0226354
R5126 VPWR VPWR.n729 0.0226354
R5127 VPWR VPWR.n762 0.0226354
R5128 VPWR VPWR.n763 0.0226354
R5129 VPWR VPWR.n785 0.0226354
R5130 VPWR VPWR.n794 0.0226354
R5131 VPWR.n830 VPWR 0.0226354
R5132 VPWR.n825 VPWR 0.0226354
R5133 VPWR.n471 VPWR 0.0226354
R5134 VPWR VPWR.n492 0.0226354
R5135 VPWR.n523 VPWR 0.0226354
R5136 VPWR VPWR.n449 0.0226354
R5137 VPWR.n674 VPWR 0.0226354
R5138 VPWR.n673 VPWR 0.0226354
R5139 VPWR.n662 VPWR 0.0226354
R5140 VPWR.n642 VPWR 0.0226354
R5141 VPWR.n635 VPWR 0.0226354
R5142 VPWR.n626 VPWR 0.0226354
R5143 VPWR VPWR.n0 0.0226354
R5144 VPWR.n1182 VPWR 0.0226354
R5145 VPWR.n1170 VPWR 0.0226354
R5146 VPWR.n1168 VPWR 0.0226354
R5147 VPWR VPWR.n137 0.0226354
R5148 VPWR.n139 VPWR 0.0226354
R5149 VPWR.n111 VPWR 0.0226354
R5150 VPWR VPWR.n183 0.0226354
R5151 VPWR VPWR.n184 0.0226354
R5152 VPWR.n285 VPWR 0.0226354
R5153 VPWR VPWR.n189 0.0226354
R5154 VPWR.n279 VPWR 0.0226354
R5155 VPWR.n274 VPWR 0.0226354
R5156 VPWR.n265 VPWR 0.0226354
R5157 VPWR.n260 VPWR 0.0226354
R5158 VPWR.n254 VPWR 0.0226354
R5159 VPWR VPWR.n73 0.0213333
R5160 VPWR VPWR.n71 0.0200312
R5161 VPWR.n874 VPWR 0.0187292
R5162 VPWR.n222 VPWR 0.0187292
R5163 VPWR.n399 VPWR.n398 0.0135208
R5164 VPWR.n371 VPWR.n31 0.0135208
R5165 VPWR.n1145 VPWR.n1144 0.0135208
R5166 VPWR.n293 VPWR.n51 0.0135208
R5167 VPWR.n1113 VPWR.n57 0.0135208
R5168 VPWR.n1097 VPWR.n71 0.0135208
R5169 VPWR.n1092 VPWR.n1077 0.0135208
R5170 VPWR.n944 VPWR.n324 0.0135208
R5171 VPWR.n320 VPWR.n317 0.0135208
R5172 VPWR.n987 VPWR.n986 0.0135208
R5173 VPWR.n99 VPWR.n96 0.0135208
R5174 VPWR.n1029 VPWR.n84 0.0135208
R5175 VPWR.n1056 VPWR.n1046 0.0135208
R5176 VPWR.n706 VPWR.n704 0.0135208
R5177 VPWR.n730 VPWR.n686 0.0135208
R5178 VPWR.n441 VPWR.n438 0.0135208
R5179 VPWR.n875 VPWR.n874 0.0135208
R5180 VPWR.n865 VPWR.n784 0.0135208
R5181 VPWR.n842 VPWR.n797 0.0135208
R5182 VPWR.n831 VPWR.n830 0.0135208
R5183 VPWR.n546 VPWR.n545 0.0135208
R5184 VPWR.n538 VPWR.n537 0.0135208
R5185 VPWR.n510 VPWR.n509 0.0135208
R5186 VPWR.n681 VPWR.n680 0.0135208
R5187 VPWR.n656 VPWR.n552 0.0135208
R5188 VPWR.n649 VPWR.n575 0.0135208
R5189 VPWR.n629 VPWR.n587 0.0135208
R5190 VPWR.n619 VPWR.n618 0.0135208
R5191 VPWR.n172 VPWR.n171 0.0135208
R5192 VPWR.n1192 VPWR.n1191 0.0135208
R5193 VPWR.n1165 VPWR.n1164 0.0135208
R5194 VPWR.n137 VPWR.n122 0.0135208
R5195 VPWR.n185 VPWR.n105 0.0135208
R5196 VPWR.n197 VPWR.n196 0.0135208
R5197 VPWR.n222 VPWR.n214 0.0135208
R5198 VPWR.n247 VPWR.n246 0.0135208
R5199 VPWR VPWR.n339 0.00961458
R5200 VPWR VPWR.n31 0.00961458
R5201 VPWR VPWR.n293 0.00961458
R5202 VPWR VPWR.n890 0.00961458
R5203 VPWR VPWR.n324 0.00961458
R5204 VPWR VPWR.n84 0.00961458
R5205 VPWR VPWR.n415 0.00961458
R5206 VPWR VPWR.n686 0.00961458
R5207 VPWR.n545 VPWR 0.00961458
R5208 VPWR VPWR.n552 0.00961458
R5209 VPWR.n172 VPWR 0.00961458
R5210 VPWR.n1164 VPWR 0.00961458
R5211 VPWR.n402 VPWR 0.0083125
R5212 VPWR VPWR.n797 0.0083125
R5213 VPWR VPWR.n485 0.0083125
R5214 VPWR VPWR.n587 0.0083125
R5215 VPWR.n77 VPWR 0.00310417
R5216 VPWR.n295 VPWR 0.00180208
R5217 VPWR.n779 VPWR 0.00180208
R5218 VPWR.n5 VPWR 0.00180208
R5219 VPWR.n190 VPWR 0.00180208
R5220 _01_.n25 _01_.n1 620.708
R5221 _01_.t18 _01_.t4 395.01
R5222 _35_.B _01_.t18 320.745
R5223 _01_.n14 _01_.t15 241.536
R5224 _01_.n2 _01_.t12 241.536
R5225 _01_.n22 _01_.t17 241.536
R5226 _01_.n20 _01_.t8 241.536
R5227 _01_.n4 _01_.t21 236.18
R5228 _01_.n6 _01_.t16 236.18
R5229 _12_.X _01_.n26 216.464
R5230 _01_.n11 _01_.t7 204.656
R5231 _01_.n17 _01_.t23 201.369
R5232 _14_.B _01_.n22 174.779
R5233 _01_.n14 _01_.t9 169.237
R5234 _01_.n2 _01_.t20 169.237
R5235 _01_.n22 _01_.t10 169.237
R5236 _01_.n20 _01_.t13 169.237
R5237 _01_.n4 _01_.t14 163.881
R5238 _01_.n6 _01_.t6 163.881
R5239 _26_.A _01_.n14 156.329
R5240 _34_.A_N _01_.n3 155.685
R5241 _37_.B _01_.n2 153.877
R5242 _01_.n5 _01_.n4 153.165
R5243 _01_.n18 _01_.n17 152.827
R5244 _01_.n12 _01_.n11 152
R5245 _01_.n10 _01_.n9 152
R5246 _01_.n7 _01_.n6 152
R5247 _01_.n21 _01_.n20 152
R5248 _01_.n3 _01_.t5 142.994
R5249 _01_.n17 _01_.t22 132.282
R5250 _01_.n3 _01_.t11 126.927
R5251 _01_.n10 _01_.t19 121.109
R5252 _01_.n11 _01_.n10 40.9982
R5253 _01_.n26 _01_.t2 38.5719
R5254 _01_.n26 _01_.t3 38.5719
R5255 _01_.n23 _14_.B 35.7985
R5256 _01_.n15 _26_.A 30.089
R5257 _01_.n23 _01_.n21 29.0338
R5258 _01_.n0 _37_.B 28.9232
R5259 _01_.n1 _01_.t0 26.5955
R5260 _01_.n1 _01_.t1 26.5955
R5261 _01_.n19 _01_.n18 16.2128
R5262 _01_.n8 _01_.n7 15.0515
R5263 _01_.n13 _32_.A_N 14.0268
R5264 _01_.n0 _01_.n5 13.0777
R5265 _01_.n0 _34_.A_N 12.5975
R5266 _01_.n15 _35_.B 12.5005
R5267 _01_.n9 _32_.A_N 10.7299
R5268 _32_.A_N _01_.n12 9.6005
R5269 _01_.n25 _01_.n24 9.3005
R5270 _01_.n13 _01_.n8 8.88649
R5271 _01_.n16 _01_.n13 8.01149
R5272 _01_.n8 _01_.n0 7.95495
R5273 _01_.n16 _01_.n15 7.25891
R5274 _01_.n19 _01_.n16 5.94006
R5275 _01_.n24 _01_.n23 5.44963
R5276 _01_.n24 _01_.n19 4.5005
R5277 _01_.n5 _31_.B 3.29747
R5278 _01_.n12 _32_.A_N 3.2005
R5279 _12_.X _01_.n25 3.2005
R5280 _01_.n21 _20_.B 2.93383
R5281 _01_.n7 _25_.B 2.52171
R5282 _01_.n9 _32_.A_N 2.07109
R5283 _01_.n18 _17_.C_N 1.75534
R5284 n_d[0].n2 n_d[0].n1 647.148
R5285 n_d[0].n7 n_d[0].n4 243.627
R5286 n_d[0].n2 n_d[0].n0 194.441
R5287 n_d[0].n6 n_d[0].n5 185
R5288 n_d[0].n5 n_d[0].t4 40.0005
R5289 n_d[0].n5 n_d[0].t5 40.0005
R5290 n_d[0].n4 n_d[0].t6 40.0005
R5291 n_d[0].n4 n_d[0].t7 40.0005
R5292 n_d[0].n6 n_d[0] 30.3501
R5293 n_d[0].n0 n_d[0].t3 27.5805
R5294 n_d[0].n0 n_d[0].t0 27.5805
R5295 n_d[0].n1 n_d[0].t1 27.5805
R5296 n_d[0].n1 n_d[0].t2 27.5805
R5297 n_d[0] n_d[0].n3 19.2609
R5298 n_d[0].n3 n_d[0].n2 15.5262
R5299 n_d[0].n7 n_d[0].n6 15.262
R5300 n_d[0].n8 n_d[0] 9.00791
R5301 n_d[0].n8 n_d[0].n7 6.77697
R5302 n_d[0].n3 n_d[0] 2.70819
R5303 n_d[0] n_d[0].n8 1.73877
R5304 y_d[0].n2 y_d[0].n0 647.148
R5305 y_d[0].n7 y_d[0].n4 200.262
R5306 y_d[0].n2 y_d[0].n1 194.441
R5307 y_d[0].n6 y_d[0].n5 185
R5308 y_d[0].n7 y_d[0].n6 58.6278
R5309 y_d[0].n5 y_d[0].t5 40.0005
R5310 y_d[0].n5 y_d[0].t6 40.0005
R5311 y_d[0].n4 y_d[0].t7 40.0005
R5312 y_d[0].n4 y_d[0].t4 40.0005
R5313 y_d[0].n1 y_d[0].t3 27.5805
R5314 y_d[0].n1 y_d[0].t0 27.5805
R5315 y_d[0].n0 y_d[0].t1 27.5805
R5316 y_d[0].n0 y_d[0].t2 27.5805
R5317 y_d[0].n6 y_d[0] 23.1558
R5318 y_d[0] y_d[0].n3 19.2609
R5319 y_d[0].n3 y_d[0].n2 15.5262
R5320 y_d[0].n8 y_d[0] 9.00791
R5321 y_d[0].n8 y_d[0].n7 6.77697
R5322 y_d[0].n3 y_d[0] 2.70819
R5323 y_d[0] y_d[0].n8 1.73877
R5324 y_d[6].n6 y_d[6].n5 647.148
R5325 y_d[6].n2 y_d[6].n0 243.627
R5326 y_d[6].n2 y_d[6].n1 200.262
R5327 y_d[6].n6 y_d[6].n4 194.441
R5328 y_d[6].n0 y_d[6].t5 40.0005
R5329 y_d[6].n0 y_d[6].t6 40.0005
R5330 y_d[6].n1 y_d[6].t7 40.0005
R5331 y_d[6].n1 y_d[6].t4 40.0005
R5332 y_d[6].n4 y_d[6].t3 27.5805
R5333 y_d[6].n4 y_d[6].t0 27.5805
R5334 y_d[6].n5 y_d[6].t1 27.5805
R5335 y_d[6].n5 y_d[6].t2 27.5805
R5336 y_d[6].n3 y_d[6] 24.7994
R5337 y_d[6] y_d[6].n6 9.86463
R5338 y_d[6].n3 y_d[6].n2 7.72512
R5339 y_d[6] y_d[6].n3 2.68692
R5340 n_d[1].n6 n_d[1].n5 647.148
R5341 n_d[1].n2 n_d[1].n0 243.627
R5342 n_d[1].n2 n_d[1].n1 200.262
R5343 n_d[1].n6 n_d[1].n4 194.441
R5344 n_d[1].n0 n_d[1].t5 40.0005
R5345 n_d[1].n0 n_d[1].t4 40.0005
R5346 n_d[1].n1 n_d[1].t6 40.0005
R5347 n_d[1].n1 n_d[1].t7 40.0005
R5348 n_d[1].n3 n_d[1] 27.6001
R5349 n_d[1].n4 n_d[1].t3 27.5805
R5350 n_d[1].n4 n_d[1].t2 27.5805
R5351 n_d[1].n5 n_d[1].t1 27.5805
R5352 n_d[1].n5 n_d[1].t0 27.5805
R5353 n_d[1].n3 n_d[1] 15.365
R5354 n_d[1] n_d[1].n2 10.4115
R5355 n_d[1] n_d[1].n6 9.86463
R5356 n_d[1] n_d[1].n3 4.18512
R5357 n_d[7].n5 n_d[7].n4 647.148
R5358 n_d[7].n2 n_d[7].n0 243.627
R5359 n_d[7].n2 n_d[7].n1 200.262
R5360 n_d[7].n5 n_d[7].n3 194.441
R5361 n_d[7].n0 n_d[7].t5 40.0005
R5362 n_d[7].n0 n_d[7].t6 40.0005
R5363 n_d[7].n1 n_d[7].t7 40.0005
R5364 n_d[7].n1 n_d[7].t4 40.0005
R5365 n_d[7].n3 n_d[7].t3 27.5805
R5366 n_d[7].n3 n_d[7].t0 27.5805
R5367 n_d[7].n4 n_d[7].t1 27.5805
R5368 n_d[7].n4 n_d[7].t2 27.5805
R5369 n_d[7] n_d[7].n6 14.9998
R5370 n_d[7] n_d[7].n5 9.86463
R5371 n_d[7].n6 n_d[7].n2 7.72512
R5372 n_d[7].n6 n_d[7] 2.68692
R5373 y_d[7].n6 y_d[7].n5 647.148
R5374 y_d[7].n2 y_d[7].n0 243.627
R5375 y_d[7].n2 y_d[7].n1 200.262
R5376 y_d[7].n6 y_d[7].n4 194.441
R5377 y_d[7].n0 y_d[7].t5 40.0005
R5378 y_d[7].n0 y_d[7].t6 40.0005
R5379 y_d[7].n1 y_d[7].t7 40.0005
R5380 y_d[7].n1 y_d[7].t4 40.0005
R5381 y_d[7].n4 y_d[7].t1 27.5805
R5382 y_d[7].n4 y_d[7].t2 27.5805
R5383 y_d[7].n5 y_d[7].t3 27.5805
R5384 y_d[7].n5 y_d[7].t0 27.5805
R5385 y_d[7].n7 y_d[7] 20.4081
R5386 y_d[7].n8 y_d[7] 19.2609
R5387 y_d[7].n7 y_d[7].n6 14.0492
R5388 y_d[7] y_d[7].n3 9.00791
R5389 y_d[7].n3 y_d[7].n2 6.77697
R5390 y_d[7] y_d[7].n8 2.70819
R5391 y_d[7].n3 y_d[7] 1.73877
R5392 y_d[7].n8 y_d[7].n7 1.47742
R5393 y_d[4].n2 y_d[4].n1 647.148
R5394 y_d[4].n7 y_d[4].n4 243.627
R5395 y_d[4].n2 y_d[4].n0 194.441
R5396 y_d[4].n6 y_d[4].n5 185
R5397 y_d[4].n5 y_d[4].t4 40.0005
R5398 y_d[4].n5 y_d[4].t5 40.0005
R5399 y_d[4].n4 y_d[4].t6 40.0005
R5400 y_d[4].n4 y_d[4].t7 40.0005
R5401 y_d[4].n0 y_d[4].t0 27.5805
R5402 y_d[4].n0 y_d[4].t1 27.5805
R5403 y_d[4].n1 y_d[4].t2 27.5805
R5404 y_d[4].n1 y_d[4].t3 27.5805
R5405 y_d[4] y_d[4].n3 19.2609
R5406 y_d[4].n6 y_d[4] 18.1191
R5407 y_d[4].n3 y_d[4].n2 15.5262
R5408 y_d[4].n7 y_d[4].n6 15.262
R5409 y_d[4].n8 y_d[4] 9.00791
R5410 y_d[4].n8 y_d[4].n7 6.77697
R5411 y_d[4].n3 y_d[4] 2.70819
R5412 y_d[4] y_d[4].n8 1.73877
R5413 y_d[2].n6 y_d[2].n5 647.148
R5414 y_d[2].n2 y_d[2].n0 243.627
R5415 y_d[2].n2 y_d[2].n1 200.262
R5416 y_d[2].n6 y_d[2].n4 194.441
R5417 y_d[2].n0 y_d[2].t6 40.0005
R5418 y_d[2].n0 y_d[2].t7 40.0005
R5419 y_d[2].n1 y_d[2].t4 40.0005
R5420 y_d[2].n1 y_d[2].t5 40.0005
R5421 y_d[2].n4 y_d[2].t1 27.5805
R5422 y_d[2].n4 y_d[2].t2 27.5805
R5423 y_d[2].n5 y_d[2].t3 27.5805
R5424 y_d[2].n5 y_d[2].t0 27.5805
R5425 y_d[2].n3 y_d[2] 23.3007
R5426 y_d[2] y_d[2].n6 9.86463
R5427 y_d[2].n3 y_d[2].n2 7.72512
R5428 y_d[2] y_d[2].n3 2.68692
R5429 y_d[5].n2 y_d[5].n1 647.148
R5430 y_d[5].n7 y_d[5].n5 243.627
R5431 y_d[5].n7 y_d[5].n6 200.262
R5432 y_d[5].n2 y_d[5].n0 194.441
R5433 y_d[5].n5 y_d[5].t7 40.0005
R5434 y_d[5].n5 y_d[5].t5 40.0005
R5435 y_d[5].n6 y_d[5].t6 40.0005
R5436 y_d[5].n6 y_d[5].t4 40.0005
R5437 y_d[5].n0 y_d[5].t1 27.5805
R5438 y_d[5].n0 y_d[5].t2 27.5805
R5439 y_d[5].n1 y_d[5].t3 27.5805
R5440 y_d[5].n1 y_d[5].t0 27.5805
R5441 y_d[5].n4 y_d[5] 27.551
R5442 y_d[5].n4 y_d[5].n3 16.5745
R5443 y_d[5].n3 y_d[5].n2 15.5262
R5444 y_d[5] y_d[5].n8 9.00791
R5445 y_d[5].n8 y_d[5].n7 6.77697
R5446 y_d[5].n3 y_d[5] 2.70819
R5447 y_d[5] y_d[5].n4 2.68692
R5448 y_d[5].n8 y_d[5] 1.73877
R5449 n_d[4].n6 n_d[4].n5 647.148
R5450 n_d[4].n3 n_d[4].n0 200.262
R5451 n_d[4].n6 n_d[4].n4 194.441
R5452 n_d[4].n2 n_d[4].n1 185
R5453 n_d[4].n3 n_d[4].n2 58.6278
R5454 n_d[4].n1 n_d[4].t4 40.0005
R5455 n_d[4].n1 n_d[4].t5 40.0005
R5456 n_d[4].n0 n_d[4].t6 40.0005
R5457 n_d[4].n0 n_d[4].t7 40.0005
R5458 n_d[4].n4 n_d[4].t2 27.5805
R5459 n_d[4].n4 n_d[4].t3 27.5805
R5460 n_d[4].n5 n_d[4].t0 27.5805
R5461 n_d[4].n5 n_d[4].t1 27.5805
R5462 n_d[4].n2 n_d[4] 19.3412
R5463 n_d[4] n_d[4].n3 10.4115
R5464 n_d[4] n_d[4].n6 9.86463
R5465 n_d[5].n6 n_d[5].n5 647.148
R5466 n_d[5].n3 n_d[5].n0 200.262
R5467 n_d[5].n6 n_d[5].n4 194.441
R5468 n_d[5].n2 n_d[5].n1 185
R5469 n_d[5].n3 n_d[5].n2 58.6278
R5470 n_d[5].n1 n_d[5].t6 40.0005
R5471 n_d[5].n1 n_d[5].t7 40.0005
R5472 n_d[5].n0 n_d[5].t4 40.0005
R5473 n_d[5].n0 n_d[5].t5 40.0005
R5474 n_d[5].n4 n_d[5].t3 27.5805
R5475 n_d[5].n4 n_d[5].t0 27.5805
R5476 n_d[5].n5 n_d[5].t1 27.5805
R5477 n_d[5].n5 n_d[5].t2 27.5805
R5478 n_d[5].n2 n_d[5] 23.7122
R5479 n_d[5] n_d[5].n3 10.4115
R5480 n_d[5] n_d[5].n6 9.86463
R5481 n_d[2].n6 n_d[2].n5 647.148
R5482 n_d[2].n3 n_d[2].n0 243.627
R5483 n_d[2].n6 n_d[2].n4 194.441
R5484 n_d[2].n2 n_d[2].n1 185
R5485 n_d[2].n1 n_d[2].t4 40.0005
R5486 n_d[2].n1 n_d[2].t7 40.0005
R5487 n_d[2].n0 n_d[2].t5 40.0005
R5488 n_d[2].n0 n_d[2].t6 40.0005
R5489 n_d[2].n4 n_d[2].t1 27.5805
R5490 n_d[2].n4 n_d[2].t3 27.5805
R5491 n_d[2].n5 n_d[2].t2 27.5805
R5492 n_d[2].n5 n_d[2].t0 27.5805
R5493 n_d[2].n2 n_d[2] 19.3412
R5494 n_d[2].n3 n_d[2].n2 15.262
R5495 n_d[2] n_d[2].n3 10.4115
R5496 n_d[2] n_d[2].n6 9.86463
R5497 y_d[3].n5 y_d[3].n4 647.148
R5498 y_d[3].n2 y_d[3].n0 243.627
R5499 y_d[3].n2 y_d[3].n1 200.262
R5500 y_d[3].n5 y_d[3].n3 194.441
R5501 y_d[3].n0 y_d[3].t6 40.0005
R5502 y_d[3].n0 y_d[3].t7 40.0005
R5503 y_d[3].n1 y_d[3].t4 40.0005
R5504 y_d[3].n1 y_d[3].t5 40.0005
R5505 y_d[3].n3 y_d[3].t1 27.5805
R5506 y_d[3].n3 y_d[3].t2 27.5805
R5507 y_d[3].n4 y_d[3].t3 27.5805
R5508 y_d[3].n4 y_d[3].t0 27.5805
R5509 y_d[3].n7 y_d[3] 22.6936
R5510 y_d[3] y_d[3].n6 19.2609
R5511 y_d[3].n6 y_d[3].n5 15.5262
R5512 y_d[3].n7 y_d[3] 8.05976
R5513 y_d[3].n8 y_d[3].n2 6.77697
R5514 y_d[3].n6 y_d[3] 2.70819
R5515 y_d[3] y_d[3].n8 1.73877
R5516 y_d[3].n8 y_d[3].n7 0.948648
R5517 y_d[1].n5 y_d[1].n4 647.148
R5518 y_d[1].n2 y_d[1].n0 243.627
R5519 y_d[1].n2 y_d[1].n1 200.262
R5520 y_d[1].n5 y_d[1].n3 194.441
R5521 y_d[1].n0 y_d[1].t6 40.0005
R5522 y_d[1].n0 y_d[1].t7 40.0005
R5523 y_d[1].n1 y_d[1].t4 40.0005
R5524 y_d[1].n1 y_d[1].t5 40.0005
R5525 y_d[1].n3 y_d[1].t1 27.5805
R5526 y_d[1].n3 y_d[1].t2 27.5805
R5527 y_d[1].n4 y_d[1].t3 27.5805
R5528 y_d[1].n4 y_d[1].t0 27.5805
R5529 y_d[1].n7 y_d[1] 22.6936
R5530 y_d[1] y_d[1].n6 19.2609
R5531 y_d[1].n6 y_d[1].n5 15.5262
R5532 y_d[1].n7 y_d[1] 8.05976
R5533 y_d[1].n8 y_d[1].n2 6.77697
R5534 y_d[1].n6 y_d[1] 2.70819
R5535 y_d[1] y_d[1].n8 1.73877
R5536 y_d[1].n8 y_d[1].n7 0.948648
R5537 n_d[6].n2 n_d[6].n0 647.148
R5538 n_d[6].n7 n_d[6].n5 243.627
R5539 n_d[6].n7 n_d[6].n6 200.262
R5540 n_d[6].n2 n_d[6].n1 194.441
R5541 n_d[6].n5 n_d[6].t6 40.0005
R5542 n_d[6].n5 n_d[6].t4 40.0005
R5543 n_d[6].n6 n_d[6].t7 40.0005
R5544 n_d[6].n6 n_d[6].t5 40.0005
R5545 n_d[6].n1 n_d[6].t3 27.5805
R5546 n_d[6].n1 n_d[6].t1 27.5805
R5547 n_d[6].n0 n_d[6].t2 27.5805
R5548 n_d[6].n0 n_d[6].t0 27.5805
R5549 n_d[6].n4 n_d[6] 20.3372
R5550 n_d[6].n4 n_d[6].n3 16.5745
R5551 n_d[6].n3 n_d[6].n2 15.5262
R5552 n_d[6] n_d[6].n8 9.00791
R5553 n_d[6].n8 n_d[6].n7 6.77697
R5554 n_d[6].n3 n_d[6] 2.70819
R5555 n_d[6] n_d[6].n4 2.68692
R5556 n_d[6].n8 n_d[6] 1.73877
R5557 in[0].n0 in[0].t0 260.322
R5558 in[0].n0 in[0].t1 175.169
R5559 in[0].n1 in[0].n0 153.385
R5560 in[0] in[0].n1 26.4102
R5561 in[0].n1 in[0] 2.94104
R5562 n_d[3].n6 n_d[3].n5 647.148
R5563 n_d[3].n2 n_d[3].n0 243.627
R5564 n_d[3].n2 n_d[3].n1 200.262
R5565 n_d[3].n6 n_d[3].n4 194.441
R5566 n_d[3].n0 n_d[3].t4 40.0005
R5567 n_d[3].n0 n_d[3].t5 40.0005
R5568 n_d[3].n1 n_d[3].t6 40.0005
R5569 n_d[3].n1 n_d[3].t7 40.0005
R5570 n_d[3].n4 n_d[3].t3 27.5805
R5571 n_d[3].n4 n_d[3].t1 27.5805
R5572 n_d[3].n5 n_d[3].t0 27.5805
R5573 n_d[3].n5 n_d[3].t2 27.5805
R5574 n_d[3].n3 n_d[3] 24.7206
R5575 n_d[3] n_d[3].n6 9.86463
R5576 n_d[3].n3 n_d[3].n2 7.72512
R5577 n_d[3] n_d[3].n3 2.68692
R5578 in[1].n0 in[1].t0 260.322
R5579 in[1].n0 in[1].t1 175.169
R5580 in[1].n1 in[1].n0 152
R5581 in[1] in[1].n1 23.2116
R5582 in[1].n1 in[1] 1.55726
R5583 in[2].n0 in[2].t0 260.322
R5584 in[2].n0 in[2].t1 175.169
R5585 in[2].n1 in[2].n0 152
R5586 in[2] in[2].n1 22.8857
R5587 in[2].n1 in[2] 1.55726
C0 _09_ _03_ 0.022129f
C1 _08_ _04_ 6.79e-20
C2 net8 a_5849_6147# 2.08e-19
C3 a_3148_4215# net15 4.51e-19
C4 a_2387_7379# a_3307_7379# 2.31e-20
C5 net17 a_4031_6740# 0.022272f
C6 a_3491_6549# _05_ 0.009119f
C7 net4 a_4307_6740# 0.115344f
C8 a_2939_6549# _03_ 2.99e-19
C9 a_2821_3561# _02_ 0.00197f
C10 _09_ net3 0.162263f
C11 a_6099_7119# _04_ 1.75e-21
C12 net13 a_2879_2223# 0.048867f
C13 a_5547_7119# net7 0.005939f
C14 net2 a_3615_4943# 0.003294f
C15 n_d[0] net17 9.58e-20
C16 net11 _03_ 3.04e-20
C17 net3 a_2939_6549# 0.011273f
C18 net2 a_4307_6740# 7.59e-20
C19 net1 a_2387_5461# 0.00906f
C20 a_3619_6147# net19 1.55e-19
C21 _02_ a_3309_5309# 0.003163f
C22 net13 net12 0.340337f
C23 net2 a_5137_2388# 0.109635f
C24 a_5547_7119# _00_ 0.001073f
C25 y_d[1] VPWR 0.419327f
C26 n_d[3] net19 3.74e-20
C27 a_2376_6263# net2 0.093667f
C28 net13 a_4167_3311# 1.43e-19
C29 a_2975_6147# _03_ 0.053532f
C30 a_5687_6740# _02_ 1.37e-19
C31 _00_ a_5476_6351# 0.002549f
C32 a_7437_2388# VPWR 0.281601f
C33 _00_ a_2869_6147# 9.44e-19
C34 y_d[7] a_2376_6263# 2.32e-19
C35 a_5297_6147# _07_ 1.99e-19
C36 VPWR a_7111_6575# 0.517103f
C37 net3 a_2975_6147# 0.320208f
C38 a_4399_7338# net5 0.131424f
C39 _04_ a_3859_7379# 0.009576f
C40 a_3289_3561# _02_ 0.002201f
C41 y_d[6] a_2376_6263# 1.65e-20
C42 _05_ net5 4.06e-19
C43 _10_ _03_ 1.46e-20
C44 _03_ net6 5.03e-19
C45 VPWR _08_ 0.198815f
C46 _09_ a_3619_6147# 0.001423f
C47 y_d[0] _00_ 6.39e-19
C48 net18 net19 0.012289f
C49 net3 net6 6.72e-19
C50 net3 _10_ 0.024506f
C51 a_6099_7119# VPWR 0.415462f
C52 _09_ n_d[3] 9.71e-21
C53 a_3701_6147# net17 2.99e-19
C54 net16 net2 0.033233f
C55 a_3384_5467# net17 1.24e-19
C56 _08_ a_3491_6549# 2.54e-19
C57 n_d[4] _04_ 4.75e-20
C58 a_3513_6147# net2 0.094679f
C59 net3 a_3342_5493# 3.24e-19
C60 net13 net2 6.97e-19
C61 net2 net9 1.82e-20
C62 n_d[7] net10 6.42e-20
C63 net8 net19 0.129236f
C64 net11 n_d[3] 4.75e-20
C65 in[0] net13 0.147979f
C66 _00_ a_2667_5175# 0.184638f
C67 net1 a_3986_5493# 4.12e-21
C68 a_6028_6351# net9 0.002837f
C69 _00_ a_2387_4373# 0.00131f
C70 a_3619_6147# a_2975_6147# 8.34e-19
C71 net3 a_3155_5056# 5.65e-19
C72 VPWR a_3859_7379# 0.414636f
C73 net18 _09_ 0.004508f
C74 _00_ a_2879_2223# 0.009027f
C75 net11 n_d[7] 0.025568f
C76 net18 a_2939_6549# 0.001138f
C77 a_3619_6147# net6 1.63e-19
C78 a_3491_6549# a_3859_7379# 0.001239f
C79 a_5849_6147# _02_ 0.105182f
C80 net8 net10 0.057549f
C81 y_d[5] _02_ 3.56e-22
C82 a_3619_6147# _10_ 6.72e-22
C83 net1 _03_ 0.115311f
C84 net12 _00_ 0.159488f
C85 n_d[3] net6 1.67e-19
C86 a_2387_7379# net2 1.47e-20
C87 a_4167_3311# _00_ 1.06e-19
C88 net3 net1 0.657665f
C89 a_2511_6147# net2 3.48e-19
C90 a_2387_7379# y_d[7] 0.021454f
C91 n_d[4] VPWR 0.458276f
C92 net16 a_3615_4943# 2.77e-20
C93 net8 net11 0.30626f
C94 a_2667_3463# VPWR 0.200835f
C95 a_2387_7379# y_d[6] 0.328904f
C96 a_3057_6147# a_2869_6147# 7.47e-21
C97 a_2387_5461# _03_ 4.34e-20
C98 y_d[2] VPWR 0.502535f
C99 a_3513_6147# a_3615_4943# 5.55e-21
C100 net17 _04_ 0.021495f
C101 n_d[1] a_3755_5639# 2.36e-22
C102 a_2667_3463# net15 3.42e-21
C103 net3 a_2387_5461# 0.004021f
C104 net18 net6 1.6e-19
C105 n_d[5] VPWR 0.44494f
C106 a_2376_6263# net16 5.95e-20
C107 a_3061_3971# a_2879_2223# 1.27e-20
C108 _02_ a_4028_5467# 0.169457f
C109 a_4031_6740# a_2387_6549# 3.78e-20
C110 net2 net7 7.05e-20
C111 a_3859_7379# net5 0.409485f
C112 a_3111_5639# a_3307_7379# 2.2e-21
C113 y_d[4] a_3755_5639# 1.75e-19
C114 a_2737_3561# VPWR 0.014462f
C115 n_d[0] a_2387_6549# 0.109428f
C116 _02_ a_5008_5487# 0.003568f
C117 _07_ _04_ 0.101419f
C118 a_4355_6147# net19 1.55e-19
C119 _02_ a_2821_4943# 0.009257f
C120 net1 a_2961_3855# 0.081244f
C121 net8 _10_ 0.052414f
C122 _00_ net2 0.301627f
C123 net8 net6 5.15e-20
C124 a_3619_6147# net1 0.155841f
C125 in[0] _00_ 9.4e-20
C126 VPWR a_3237_5309# 3.4e-20
C127 a_3755_5639# a_4028_5467# 0.167615f
C128 a_3111_5639# a_3261_5493# 0.002605f
C129 _00_ a_6028_6351# 0.001512f
C130 VPWR a_5437_6575# 1.6e-19
C131 n_d[4] net5 0.001826f
C132 a_2387_3027# _02_ 0.037144f
C133 _02_ net19 0.059371f
C134 _08_ a_3309_5309# 2.57e-19
C135 VPWR net17 0.276872f
C136 a_4355_6147# a_4437_6147# 0.004937f
C137 a_3707_3311# _02_ 0.040522f
C138 a_3019_7338# n_d[0] 8.51e-20
C139 a_2511_6147# a_2376_6263# 0.008678f
C140 a_3019_7338# n_d[2] 0.039283f
C141 a_3491_6549# net17 0.202955f
C142 in[2] net3 0.003035f
C143 net18 net1 1.54e-20
C144 a_3755_5639# net19 2.68e-22
C145 y_d[3] a_2387_5461# 8.68e-20
C146 VPWR _07_ 0.350367f
C147 y_d[5] _05_ 1.52e-19
C148 net2 a_3061_3971# 0.218627f
C149 n_d[1] a_4399_7338# 5.94e-19
C150 a_2607_6147# net1 4.44e-19
C151 a_5547_7119# a_5297_6147# 1.96e-20
C152 a_4249_6147# net2 0.102373f
C153 net10 _02_ 0.120505f
C154 net3 a_3986_5493# 5e-19
C155 a_6099_7119# a_6651_7119# 0.003298f
C156 n_d[1] _05_ 4.07e-19
C157 _09_ _02_ 1.23e-19
C158 a_5297_6147# a_5476_6351# 0.007688f
C159 _02_ a_2939_6549# 7e-20
C160 n_d[0] a_2869_6147# 4.64e-19
C161 a_4903_6575# net4 5.28e-19
C162 _00_ a_3615_4943# 0.029099f
C163 a_2667_3463# a_3219_3463# 0.001119f
C164 a_5547_7119# n_d[6] 2.31e-21
C165 net3 _03_ 0.596753f
C166 net11 _02_ 0.081905f
C167 _09_ a_3129_6147# 5.2e-19
C168 a_5560_6351# _02_ 3.2e-19
C169 _05_ a_4028_5467# 7.47e-20
C170 a_2667_3463# a_2821_3561# 0.010303f
C171 a_2975_6147# _02_ 8.99e-22
C172 n_d[2] a_3307_7379# 0.337274f
C173 a_3057_6147# net2 2.04e-19
C174 net2 a_3111_5639# 0.097352f
C175 n_d[4] a_5687_6740# 9.32e-20
C176 _02_ net6 4.24e-20
C177 _10_ _02_ 0.169021f
C178 a_3129_6147# a_2975_6147# 0.008535f
C179 y_d[5] _08_ 3.58e-19
C180 n_d[4] a_6651_7119# 2.04e-19
C181 net9 net7 1.25e-19
C182 n_d[3] a_4779_7379# 0.3328f
C183 a_4745_5533# net7 0.137606f
C184 _00_ net16 0.002429f
C185 a_3619_6147# _03_ 0.059264f
C186 a_4249_6147# a_4307_6740# 0.001457f
C187 _05_ net19 0.100007f
C188 a_3513_6147# _00_ 7.03e-22
C189 net3 a_2961_3855# 2.79e-21
C190 net13 _00_ 0.288591f
C191 a_3619_6147# net3 0.275853f
C192 _00_ a_4745_5533# 0.12395f
C193 y_d[4] _08_ 0.001932f
C194 _00_ net9 0.02542f
C195 a_3384_5467# a_3307_7379# 4.37e-19
C196 _10_ a_3755_5639# 3.51e-21
C197 n_d[3] net3 0.002257f
C198 n_d[5] a_6651_7119# 0.337855f
C199 _02_ a_3155_5056# 0.244359f
C200 net1 a_3571_4074# 0.035248f
C201 n_d[7] a_4779_7379# 3.67e-20
C202 a_4355_6147# net1 0.264989f
C203 a_4903_6575# a_4307_6740# 0.002227f
C204 VPWR a_2737_4943# 0.015007f
C205 a_3773_6147# _04_ 0.00109f
C206 y_d[1] a_2387_2197# 0.329593f
C207 y_d[3] net3 3.65e-20
C208 _09_ a_4399_7338# 5.35e-19
C209 _09_ _05_ 0.004171f
C210 VPWR a_3045_2767# 0.001585f
C211 y_d[1] a_2387_3027# 8.94e-19
C212 n_d[1] a_3859_7379# 0.339535f
C213 net17 a_3309_5309# 4.73e-20
C214 a_2939_6549# _05_ 8.97e-20
C215 net4 a_4031_6740# 0.146829f
C216 net1 _02_ 0.05595f
C217 net14 _02_ 0.034031f
C218 a_3373_3561# VPWR 0.008908f
C219 VPWR a_2387_6549# 0.454473f
C220 a_5547_7119# _04_ 1.68e-20
C221 net8 a_4779_7379# 2.84e-19
C222 a_7111_6575# net19 4.14e-20
C223 y_d[0] a_2961_2767# 1.02e-20
C224 net13 a_3061_3971# 6.1e-19
C225 net8 _03_ 1.45e-19
C226 n_d[0] net4 0.016054f
C227 net11 _05_ 1.98e-20
C228 a_2607_6147# net3 0.00267f
C229 net2 a_4031_6740# 0.001165f
C230 a_4443_3855# net2 0.038895f
C231 a_2869_6147# _04_ 5.29e-20
C232 _08_ net19 2.07e-20
C233 n_d[2] net4 2.52e-19
C234 y_d[7] a_4031_6740# 6.98e-20
C235 a_4028_5467# a_3859_7379# 1.85e-21
C236 n_d[1] n_d[4] 1.79e-21
C237 net2 _06_ 0.208301f
C238 a_3129_6147# net1 8.41e-19
C239 a_2975_6147# _05_ 2.06e-19
C240 n_d[0] net2 0.003331f
C241 a_3707_3311# _08_ 1.35e-19
C242 a_2387_5461# _02_ 0.002062f
C243 net1 a_3755_5639# 0.079733f
C244 VPWR a_3773_6147# 2.63e-19
C245 n_d[2] net2 2.79e-19
C246 y_d[7] n_d[0] 0.143217f
C247 _04_ a_3307_7379# 8.75e-19
C248 a_4399_7338# net6 0.001017f
C249 a_3019_7338# VPWR 0.242915f
C250 _00_ net7 0.157409f
C251 net10 a_7111_6575# 0.226294f
C252 n_d[2] y_d[7] 0.313736f
C253 n_d[3] n_d[7] 4.34e-20
C254 y_d[6] n_d[0] 0.1964f
C255 _05_ net6 0.022873f
C256 net16 a_3111_5639# 0.008905f
C257 y_d[6] n_d[2] 1.73e-20
C258 _09_ _08_ 1.66e-19
C259 net18 n_d[3] 3.91e-22
C260 a_5547_7119# VPWR 0.53318f
C261 net11 a_7111_6575# 2.2e-19
C262 net19 a_3859_7379# 6.23e-20
C263 a_3384_5467# net4 1.56e-20
C264 net12 a_2961_2767# 0.012296f
C265 VPWR a_5476_6351# 3.83e-19
C266 VPWR a_2869_6147# 0.09278f
C267 net8 n_d[3] 1.2e-19
C268 net2 a_3384_5467# 0.090636f
C269 a_4031_6740# a_4307_6740# 5.07e-19
C270 y_d[5] net17 0.023893f
C271 net11 a_6099_7119# 0.228016f
C272 n_d[1] net17 9.01e-19
C273 VPWR a_3307_7379# 0.417167f
C274 a_2667_3463# a_2387_2197# 1.66e-20
C275 y_d[0] VPWR 0.359804f
C276 y_d[2] a_2387_2197# 8.94e-19
C277 n_d[0] a_4307_6740# 9.96e-21
C278 a_4355_6147# _03_ 0.035636f
C279 _10_ a_7111_6575# 1.33e-19
C280 net8 n_d[7] 7.02e-20
C281 net1 a_4399_7338# 1.2e-20
C282 a_3019_7338# net5 1.36e-19
C283 _09_ a_3859_7379# 5.66e-20
C284 _00_ a_3061_3971# 0.036522f
C285 _02_ a_3986_5493# 8.98e-20
C286 a_3219_3463# a_3373_3561# 0.010303f
C287 a_2667_3463# a_2387_3027# 7.14e-19
C288 y_d[2] a_2387_3027# 0.329274f
C289 y_d[4] net17 2.61e-20
C290 net3 a_3571_4074# 5.66e-20
C291 a_3491_6549# a_3307_7379# 0.017402f
C292 net1 _05_ 0.027624f
C293 a_4355_6147# net3 0.03947f
C294 VPWR a_3261_5493# 2.46e-19
C295 n_d[0] a_2376_6263# 1.77e-20
C296 _08_ net6 1.19e-20
C297 _10_ _08_ 0.042943f
C298 a_4903_6575# net7 0.012104f
C299 a_5547_7119# net5 1.59e-20
C300 _02_ _03_ 1.51e-19
C301 VPWR a_2667_5175# 0.216131f
C302 _08_ a_3342_5493# 1.23e-19
C303 a_3755_5639# a_3986_5493# 0.004898f
C304 a_4509_6147# _04_ 0.001514f
C305 VPWR a_2387_4373# 0.532617f
C306 _00_ a_4903_6575# 2.72e-19
C307 net15 a_2667_5175# 0.001285f
C308 net15 a_2387_4373# 0.2262f
C309 net3 _02_ 0.341653f
C310 VPWR a_2879_2223# 0.379525f
C311 net4 _04_ 0.004865f
C312 _08_ a_3155_5056# 0.026979f
C313 y_d[1] net1 9.01e-20
C314 n_d[5] net10 4.97e-20
C315 n_d[0] net16 1.66e-21
C316 a_3755_5639# _03_ 3.35e-21
C317 net11 n_d[4] 0.008049f
C318 net12 VPWR 0.412615f
C319 a_2961_3855# a_3571_4074# 2.28e-20
C320 net2 _04_ 0.289566f
C321 a_3307_7379# net5 0.00101f
C322 a_5437_6575# net19 0.001078f
C323 net6 a_3859_7379# 0.03111f
C324 _00_ a_3111_5639# 0.002116f
C325 a_4167_3311# VPWR 0.325153f
C326 a_3129_6147# net3 0.004045f
C327 a_3619_6147# a_4355_6147# 7.25e-19
C328 net3 a_3755_5639# 0.262138f
C329 a_3220_4215# net2 0.004863f
C330 n_d[3] a_4355_6147# 1.26e-19
C331 y_d[7] _04_ 3.97e-20
C332 net17 net19 0.066786f
C333 net11 n_d[5] 1.97e-19
C334 net1 _08_ 0.038099f
C335 _02_ a_2961_3855# 0.016216f
C336 VPWR a_4509_6147# 2.4e-19
C337 a_3619_6147# _02_ 9.62e-22
C338 n_d[6] net9 0.039885f
C339 n_d[4] _10_ 4.03e-19
C340 _07_ net19 0.102218f
C341 VPWR net4 0.331113f
C342 a_3219_3463# y_d[0] 1.48e-19
C343 a_2387_7379# n_d[0] 2.62e-20
C344 net16 a_3384_5467# 2.71e-20
C345 a_2387_5461# _08_ 1.92e-19
C346 _09_ net17 0.02551f
C347 y_d[3] _02_ 0.008434f
C348 a_2387_7379# n_d[2] 5.46e-20
C349 VPWR net2 3.35419f
C350 a_3701_6147# a_3513_6147# 7.47e-21
C351 a_2939_6549# net17 8.47e-19
C352 net4 a_3491_6549# 0.121037f
C353 net11 a_5437_6575# 0.011723f
C354 a_3619_6147# a_3755_5639# 3.1e-20
C355 a_5547_7119# a_5687_6740# 0.010769f
C356 in[0] VPWR 0.562802f
C357 VPWR a_6028_6351# 7.61e-19
C358 net2 net15 0.367103f
C359 a_4399_7338# a_4779_7379# 3.18e-19
C360 net1 a_3859_7379# 2.89e-19
C361 y_d[7] VPWR 0.793311f
C362 net11 net17 2.75e-21
C363 net2 a_3491_6549# 0.004036f
C364 a_4307_6740# _04_ 0.00912f
C365 _03_ a_4399_7338# 0.011898f
C366 y_d[6] VPWR 0.418911f
C367 _05_ _03_ 0.107536f
C368 y_d[7] a_3491_6549# 1.77e-19
C369 y_d[5] a_2387_6549# 0.054072f
C370 a_2975_6147# net17 0.001052f
C371 a_5297_6147# net7 0.004018f
C372 a_3219_3463# a_2879_2223# 0.001294f
C373 a_4443_3855# _00_ 0.174506f
C374 n_d[1] a_2387_6549# 1.01e-19
C375 in[2] a_7437_2388# 0.195629f
C376 net3 _05_ 0.018016f
C377 net11 _07_ 2.73e-19
C378 net8 _02_ 0.056023f
C379 _00_ _06_ 0.011673f
C380 n_d[0] _00_ 7.18e-21
C381 a_5297_6147# _00_ 0.093344f
C382 net4 net5 1.93e-19
C383 net17 net6 0.008537f
C384 net13 a_2961_2767# 2.43e-19
C385 VPWR a_3905_5493# 1.59e-19
C386 y_d[4] a_2387_6549# 0.001012f
C387 _10_ net17 0.021624f
C388 a_2667_3463# net14 0.150649f
C389 y_d[2] net14 0.042113f
C390 a_2667_3463# net1 1.47e-19
C391 a_3155_5056# a_3237_5309# 0.005167f
C392 net2 net5 1.98e-21
C393 net17 a_3342_5493# 7.01e-21
C394 VPWR a_3615_4943# 0.189789f
C395 _07_ net6 4.58e-20
C396 a_3019_7338# n_d[1] 0.044512f
C397 VPWR a_4307_6740# 0.259026f
C398 y_d[7] net5 1.74e-19
C399 net14 a_2737_3561# 0.00346f
C400 a_3513_6147# _04_ 0.020587f
C401 VPWR a_5137_2388# 0.253289f
C402 net17 a_3155_5056# 4.31e-19
C403 a_3491_6549# a_3615_4943# 2.27e-20
C404 n_d[3] a_4399_7338# 0.012777f
C405 a_2376_6263# VPWR 0.197704f
C406 net3 a_7437_2388# 0.11065f
C407 a_5547_7119# a_5849_6147# 6.11e-20
C408 a_3148_4215# a_2961_3855# 1.84e-19
C409 a_3619_6147# _05_ 0.102485f
C410 _08_ _03_ 3.74e-20
C411 a_3061_3971# _06_ 0.112825f
C412 a_2387_3027# a_3045_2767# 4.66e-20
C413 a_5547_7119# n_d[1] 5.95e-22
C414 _00_ a_3384_5467# 3.11e-20
C415 net3 _08_ 0.100455f
C416 a_3219_3463# net2 0.002444f
C417 a_3219_3463# in[0] 1.04e-21
C418 a_2387_6549# net19 0.208337f
C419 net1 net17 0.437005f
C420 a_3373_3561# a_3707_3311# 3.88e-19
C421 y_d[5] a_3307_7379# 0.001317f
C422 VPWR net16 0.414648f
C423 _02_ a_3571_4074# 5.03e-20
C424 a_4355_6147# _02_ 2e-19
C425 a_4779_7379# a_3859_7379# 2.31e-20
C426 n_d[1] a_3307_7379# 0.167145f
C427 a_3513_6147# VPWR 0.086139f
C428 net16 net15 0.001073f
C429 _03_ a_3859_7379# 3.05e-20
C430 a_4307_6740# net5 3.35e-19
C431 net13 VPWR 0.315732f
C432 net1 _07_ 0.002892f
C433 VPWR net9 0.836328f
C434 VPWR a_4745_5533# 0.205805f
C435 in[1] net2 0.008337f
C436 net2 a_3309_5309# 4.11e-19
C437 net3 a_3859_7379# 4.97e-20
C438 _09_ a_2387_6549# 0.003348f
C439 net13 net15 0.00412f
C440 a_3513_6147# a_3491_6549# 0.011876f
C441 n_d[0] a_3111_5639# 7.35e-21
C442 a_3619_6147# _08_ 1.14e-19
C443 a_2939_6549# a_2387_6549# 0.003298f
C444 n_d[4] a_4779_7379# 0.001762f
C445 _04_ net7 0.055645f
C446 y_d[4] a_3261_5493# 1.93e-19
C447 n_d[7] a_7111_6575# 4.03e-20
C448 a_3289_3561# net2 4.47e-20
C449 a_6099_7119# n_d[3] 5.68e-20
C450 a_2387_7379# VPWR 0.412323f
C451 y_d[4] a_2387_4373# 0.002087f
C452 a_3755_5639# _02_ 0.01899f
C453 _10_ a_4924_5487# 2.32e-19
C454 a_2869_6147# net19 1.1e-20
C455 a_3019_7338# _09_ 0.1931f
C456 a_2511_6147# VPWR 0.001075f
C457 a_3220_4215# _00_ 2.42e-20
C458 y_d[0] a_2387_2197# 0.007264f
C459 a_3019_7338# a_2939_6549# 0.011678f
C460 a_6099_7119# n_d[7] 0.328945f
C461 a_3619_6147# a_3859_7379# 0.001184f
C462 a_5547_7119# net10 2.77e-19
C463 net8 a_7111_6575# 1.5e-19
C464 net19 a_3307_7379# 5.37e-20
C465 a_2387_6549# net6 2.63e-19
C466 y_d[0] a_2387_3027# 1.03e-19
C467 n_d[3] a_3859_7379# 0.002245f
C468 a_3111_5639# a_3384_5467# 0.167615f
C469 a_5476_6351# net10 0.001923f
C470 a_2667_5175# a_2821_4943# 0.010303f
C471 VPWR net7 0.853667f
C472 _09_ a_2869_6147# 6.16e-19
C473 in[1] a_5137_2388# 0.221617f
C474 y_d[5] net4 0.259724f
C475 net8 a_6099_7119# 0.006936f
C476 a_5547_7119# net11 0.023056f
C477 a_2869_6147# a_2939_6549# 0.012653f
C478 a_4249_6147# _04_ 0.013323f
C479 _00_ VPWR 1.98913f
C480 n_d[1] net4 6.72e-21
C481 a_2387_2197# a_2879_2223# 0.18179f
C482 _00_ a_5353_6575# 2.54e-19
C483 n_d[3] n_d[4] 0.126574f
C484 n_d[0] a_4031_6740# 4.59e-20
C485 a_2667_3463# a_2961_3855# 2.67e-19
C486 a_4443_3855# _06_ 4.32e-19
C487 a_3220_4215# a_3061_3971# 0.002605f
C488 y_d[5] net2 0.001391f
C489 a_4355_6147# _05_ 0.001196f
C490 a_3019_7338# net6 1.14e-19
C491 net17 _03_ 0.031661f
C492 a_2387_7379# net5 2.82e-21
C493 net18 a_3859_7379# 1.22e-19
C494 _09_ a_3307_7379# 0.032162f
C495 _00_ net15 0.182308f
C496 a_3219_3463# net13 0.142278f
C497 a_2939_6549# a_3307_7379# 0.001239f
C498 a_5849_6147# a_6028_6351# 0.007688f
C499 n_d[1] net2 2.04e-19
C500 _00_ a_3491_6549# 3.91e-21
C501 net12 a_2387_2197# 0.011305f
C502 y_d[7] y_d[5] 0.361483f
C503 net3 net17 0.213037f
C504 a_2869_6147# a_2975_6147# 0.13675f
C505 _07_ a_4779_7379# 0.012239f
C506 a_4903_6575# _04_ 0.003352f
C507 a_2387_3027# net12 0.120337f
C508 n_d[4] n_d[7] 0.00103f
C509 y_d[6] y_d[5] 0.10387f
C510 n_d[1] y_d[7] 0.149492f
C511 y_d[4] net2 0.001971f
C512 a_5547_7119# _10_ 0.012522f
C513 _07_ _03_ 0.023582f
C514 y_d[3] y_d[2] 0.114081f
C515 _02_ _05_ 4.33e-20
C516 net4 a_4028_5467# 2.65e-21
C517 net13 a_2821_3561# 3.88e-19
C518 y_d[6] n_d[1] 0.241626f
C519 a_3373_3561# net1 0.001168f
C520 net1 a_2387_6549# 0.010573f
C521 net16 a_3309_5309# 3.13e-20
C522 y_d[7] y_d[4] 0.001551f
C523 a_3707_3311# a_4167_3311# 0.001607f
C524 net3 _07_ 0.00931f
C525 net2 a_4028_5467# 4.11e-19
C526 a_2939_6549# a_2667_5175# 1.54e-20
C527 a_3057_6147# _04_ 7.03e-20
C528 net7 net5 9.47e-20
C529 n_d[7] n_d[5] 0.112125f
C530 y_d[6] y_d[4] 7.02e-20
C531 VPWR a_3061_3971# 0.2216f
C532 a_4249_6147# VPWR 0.101518f
C533 a_2387_5461# a_2387_6549# 0.001583f
C534 net15 a_3061_3971# 0.032637f
C535 net8 n_d[4] 0.129018f
C536 a_3307_7379# net6 0.223504f
C537 a_5687_6740# net9 4.02e-20
C538 net1 a_3773_6147# 6.08e-19
C539 a_3619_6147# net17 0.016769f
C540 _08_ a_3571_4074# 4.16e-19
C541 net4 net19 0.285122f
C542 y_d[5] a_3615_4943# 4.67e-22
C543 net13 a_3289_3561# 0.003264f
C544 net9 a_6651_7119# 0.227856f
C545 in[0] a_2387_2197# 0.088701f
C546 VPWR a_4903_6575# 0.243068f
C547 y_d[4] a_3905_5493# 3.31e-20
C548 n_d[2] a_3384_5467# 6.02e-21
C549 net8 n_d[5] 3.69e-20
C550 net2 net19 0.004237f
C551 in[0] a_2387_3027# 1.01e-19
C552 a_3707_3311# net2 0.015566f
C553 _10_ a_2667_5175# 4.05e-19
C554 _08_ _02_ 0.122114f
C555 y_d[7] net19 0.029921f
C556 n_d[3] _07_ 9.01e-19
C557 n_d[1] a_2376_6263# 4.63e-22
C558 a_3057_6147# VPWR 1.16e-19
C559 VPWR a_3111_5639# 0.206134f
C560 a_3219_3463# _00_ 0.054461f
C561 y_d[0] a_3431_2223# 0.028767f
C562 net1 a_2869_6147# 0.094612f
C563 _09_ net4 0.012562f
C564 y_d[4] a_2376_6263# 0.003485f
C565 a_2939_6549# net4 0.212039f
C566 a_4249_6147# net5 1.1e-19
C567 net8 a_5437_6575# 6.15e-20
C568 a_4437_6147# net2 2.01e-19
C569 net2 net10 9.8e-20
C570 _09_ net2 0.29681f
C571 a_3755_5639# _08_ 0.088996f
C572 a_2821_3561# _00_ 0.001572f
C573 net1 a_3307_7379# 9.82e-21
C574 a_2667_5175# a_3155_5056# 0.062241f
C575 y_d[0] net1 0.001211f
C576 a_6028_6351# net10 7.04e-19
C577 net11 net4 3.52e-20
C578 net8 net17 2.73e-20
C579 net2 a_2939_6549# 0.012647f
C580 a_4031_6740# _04_ 0.002848f
C581 _09_ y_d[7] 0.149255f
C582 y_d[5] a_3513_6147# 3e-19
C583 a_5687_6740# net7 0.001616f
C584 _02_ a_3859_7379# 4.88e-20
C585 y_d[7] a_2939_6549# 0.012794f
C586 _00_ a_3309_5309# 1.1e-19
C587 a_5849_6147# net9 0.137671f
C588 n_d[0] _04_ 2.14e-20
C589 _09_ y_d[6] 1.13e-19
C590 net3 a_4924_5487# 5.23e-19
C591 a_2975_6147# net4 0.011988f
C592 a_2879_2223# a_3431_2223# 0.001868f
C593 y_d[4] net16 0.044291f
C594 _00_ a_5687_6740# 0.025483f
C595 net8 _07_ 0.004062f
C596 a_3219_3463# a_3061_3971# 5.92e-19
C597 n_d[2] _04_ 2.2e-20
C598 net2 a_2975_6147# 0.181408f
C599 net1 a_2667_5175# 6.52e-20
C600 _03_ a_2387_6549# 1.84e-19
C601 a_4307_6740# net19 0.033296f
C602 net1 a_2387_4373# 1.36e-21
C603 net14 a_2387_4373# 1.19e-21
C604 net4 net6 0.143949f
C605 net12 a_3431_2223# 1.65e-20
C606 a_3289_3561# _00_ 0.001825f
C607 a_3755_5639# a_3859_7379# 1.92e-20
C608 net3 a_2387_6549# 0.010176f
C609 a_2376_6263# net19 1.49e-19
C610 net16 a_4028_5467# 1.67e-21
C611 y_d[7] a_2975_6147# 7.27e-19
C612 n_d[4] _02_ 9.7e-20
C613 net1 a_2879_2223# 0.001624f
C614 net2 net6 1.05e-20
C615 net2 _10_ 0.0061f
C616 net12 net14 0.003618f
C617 a_2387_5461# a_2667_5175# 7.14e-19
C618 a_4745_5533# a_4028_5467# 1.01e-19
C619 net12 net1 2.28e-19
C620 a_2667_3463# _02_ 0.132972f
C621 a_2387_5461# a_2387_4373# 0.002813f
C622 y_d[2] _02_ 2.56e-19
C623 net16 a_2821_4943# 0.002266f
C624 VPWR a_4031_6740# 0.216638f
C625 a_6028_6351# _10_ 0.001113f
C626 a_2387_7379# n_d[1] 0.092512f
C627 y_d[7] net6 5.31e-19
C628 a_4167_3311# net1 0.002202f
C629 a_4443_3855# VPWR 0.318955f
C630 _09_ a_4307_6740# 3.91e-19
C631 net2 a_3342_5493# 1.78e-19
C632 a_3701_6147# _04_ 6.12e-19
C633 a_3384_5467# _04_ 1.21e-19
C634 VPWR _06_ 0.213942f
C635 a_2387_7379# y_d[4] 4.44e-20
C636 a_4745_5533# a_5008_5487# 0.010598f
C637 a_4443_3855# net15 1.22e-19
C638 n_d[0] VPWR 0.35591f
C639 a_5297_6147# VPWR 0.172617f
C640 net3 a_3773_6147# 0.003136f
C641 a_3491_6549# a_4031_6740# 0.003294f
C642 a_2737_3561# _02_ 0.001402f
C643 a_3019_7338# net3 2.85e-19
C644 _09_ a_2376_6263# 3.14e-19
C645 net13 a_2387_2197# 0.216582f
C646 net16 net19 0.001076f
C647 net15 _06_ 0.226529f
C648 n_d[2] VPWR 0.380649f
C649 net2 a_3155_5056# 0.023253f
C650 n_d[0] a_3491_6549# 9.83e-20
C651 net11 a_4307_6740# 7.49e-20
C652 net1 a_4509_6147# 0.002917f
C653 a_4355_6147# net17 2.04e-19
C654 a_3513_6147# net19 3.41e-20
C655 net2 a_3431_2223# 4.11e-21
C656 _02_ a_3237_5309# 0.001597f
C657 net13 a_2387_3027# 4.49e-19
C658 n_d[6] VPWR 0.686834f
C659 net9 net19 1.69e-20
C660 in[0] a_3431_2223# 0.205512f
C661 a_4745_5533# net19 5.87e-21
C662 n_d[2] a_3491_6549# 6.95e-19
C663 net1 net4 7.52e-20
C664 a_2869_6147# _03_ 0.030887f
C665 net13 a_3707_3311# 0.002502f
C666 n_d[1] net7 1.98e-20
C667 a_5437_6575# _02_ 1.67e-19
C668 a_5687_6740# a_4903_6575# 0.001761f
C669 _00_ a_5849_6147# 0.078044f
C670 a_4355_6147# _07_ 0.102593f
C671 a_2376_6263# a_2975_6147# 5.82e-19
C672 net3 a_2869_6147# 0.059202f
C673 _02_ net17 0.065146f
C674 net1 net2 1.03327f
C675 a_4399_7338# a_3859_7379# 0.003294f
C676 in[0] net1 0.003451f
C677 in[0] net14 7.59e-21
C678 _10_ a_3615_4943# 0.127937f
C679 _09_ net16 0.002681f
C680 _05_ a_3859_7379# 0.010141f
C681 a_4031_6740# net5 1.73e-20
C682 a_4307_6740# net6 7.64e-19
C683 _03_ a_3307_7379# 2.96e-20
C684 a_3619_6147# a_3773_6147# 0.008535f
C685 a_3701_6147# VPWR 1.61e-19
C686 y_d[7] net1 3.52e-19
C687 VPWR a_3384_5467# 0.166515f
C688 net10 net9 0.037093f
C689 _09_ a_3513_6147# 0.001512f
C690 a_2387_7379# net19 1.11e-19
C691 a_4028_5467# net7 9.98e-20
C692 net3 a_3307_7379# 1.45e-20
C693 net18 a_2387_6549# 1.11e-19
C694 a_3019_7338# n_d[3] 4.1e-20
C695 a_2387_5461# net2 0.008513f
C696 _07_ _02_ 0.00125f
C697 a_3384_5467# a_3491_6549# 1.42e-19
C698 a_3755_5639# net17 0.013743f
C699 n_d[2] net5 0.003167f
C700 n_d[4] a_4399_7338# 1.05e-19
C701 _00_ a_4028_5467# 1.4e-19
C702 a_5008_5487# net7 0.00411f
C703 y_d[7] a_2387_5461# 8.2e-20
C704 net3 a_3261_5493# 0.005326f
C705 net11 net9 0.046616f
C706 a_5547_7119# n_d[3] 2.33e-19
C707 _00_ a_5008_5487# 0.001217f
C708 a_3513_6147# a_2975_6147# 0.001036f
C709 net1 a_3905_5493# 5.19e-19
C710 net3 a_2667_5175# 2.59e-19
C711 net18 a_3019_7338# 0.127919f
C712 VPWR a_2961_2767# 0.002283f
C713 a_2387_7379# _09_ 0.001082f
C714 net19 net7 0.023885f
C715 a_3431_2223# a_5137_2388# 2.29e-19
C716 net16 _10_ 2.33e-20
C717 a_5547_7119# n_d[7] 1.39e-19
C718 y_d[0] a_2961_3855# 1.7e-20
C719 net1 a_3615_4943# 0.005953f
C720 a_3513_6147# net6 3.13e-20
C721 a_3513_6147# _10_ 6.19e-22
C722 _00_ net19 0.081779f
C723 a_2387_3027# _00_ 6.61e-19
C724 net1 a_4307_6740# 6.56e-20
C725 n_d[3] a_3307_7379# 6.59e-19
C726 _10_ net9 0.031889f
C727 _10_ a_4745_5533# 3.02e-19
C728 net1 a_5137_2388# 4.11e-21
C729 a_3707_3311# _00_ 0.001981f
C730 a_2376_6263# net1 0.144619f
C731 VPWR _04_ 0.69792f
C732 y_d[1] y_d[2] 0.11727f
C733 net16 a_3155_5056# 4.93e-19
C734 net8 a_5547_7119# 0.272184f
C735 a_3220_4215# VPWR 2.24e-19
C736 a_2607_6147# a_2869_6147# 5.23e-21
C737 a_3491_6549# _04_ 0.001882f
C738 _00_ net10 0.188756f
C739 a_3220_4215# net15 0.002179f
C740 net18 a_3307_7379# 0.001239f
C741 net17 _05_ 0.087752f
C742 net3 a_4509_6147# 8.99e-19
C743 _09_ _00_ 0.00407f
C744 a_2376_6263# a_2387_5461# 0.010596f
C745 net4 _03_ 0.005453f
C746 a_2961_3855# a_2879_2223# 1.02e-21
C747 a_5297_6147# a_5687_6740# 0.001028f
C748 a_6099_7119# n_d[4] 0.079007f
C749 net11 net7 0.009487f
C750 net13 a_3431_2223# 0.006182f
C751 _00_ a_2939_6549# 1.58e-19
C752 y_d[4] a_3111_5639# 9.62e-19
C753 net3 net4 1.06e-19
C754 net12 a_2961_3855# 8.45e-20
C755 y_d[3] a_2387_4373# 0.32983f
C756 net1 net16 3.1e-19
C757 net2 _03_ 0.675804f
C758 _02_ a_4924_5487# 0.002639f
C759 a_4249_6147# net19 1.51e-19
C760 _02_ a_2737_4943# 0.00374f
C761 net11 _00_ 0.107906f
C762 a_3513_6147# net1 0.10031f
C763 _07_ _05_ 0.003185f
C764 y_d[7] _03_ 1.15e-19
C765 net3 net2 1.0792f
C766 a_6099_7119# n_d[5] 0.001819f
C767 net13 net1 0.063726f
C768 net13 net14 0.019852f
C769 net1 a_4745_5533# 2.99e-20
C770 _00_ a_5560_6351# 0.00592f
C771 _00_ a_2975_6147# 1.19e-19
C772 VPWR a_5353_6575# 2.56e-19
C773 y_d[7] net3 0.003299f
C774 n_d[6] a_6651_7119# 0.005112f
C775 a_2387_5461# net16 0.2073f
C776 net7 net6 1.16e-20
C777 n_d[4] a_3859_7379# 8.99e-21
C778 _04_ net5 0.009669f
C779 a_4903_6575# net19 0.033722f
C780 a_3373_3561# _02_ 0.003236f
C781 VPWR net15 0.326349f
C782 _10_ net7 0.00127f
C783 y_d[6] net3 1.65e-19
C784 a_4249_6147# a_4437_6147# 7.47e-21
C785 VPWR a_3491_6549# 0.354271f
C786 _00_ net6 1.63e-20
C787 _00_ _10_ 0.737416f
C788 a_3619_6147# net4 6.49e-20
C789 a_2387_7379# net1 1.73e-19
C790 _08_ net17 0.131764f
C791 a_3111_5639# net19 2.35e-22
C792 net2 a_2961_3855# 0.001878f
C793 y_d[5] a_4031_6740# 1.27e-19
C794 in[0] a_2961_3855# 9.87e-22
C795 a_2511_6147# net1 4.89e-19
C796 a_3619_6147# net2 0.026767f
C797 net3 a_3905_5493# 0.005328f
C798 a_3615_4943# _03_ 1.71e-22
C799 n_d[1] a_4031_6740# 2.26e-19
C800 n_d[0] y_d[5] 0.5105f
C801 a_5297_6147# a_5849_6147# 0.001113f
C802 a_4307_6740# _03_ 0.194036f
C803 _00_ a_3155_5056# 0.264455f
C804 a_6112_6351# net9 0.005795f
C805 net3 a_3615_4943# 4.96e-19
C806 n_d[1] n_d[0] 0.098807f
C807 n_d[4] n_d[5] 0.096452f
C808 VPWR net5 0.239168f
C809 a_2667_3463# y_d[2] 4.86e-21
C810 net3 a_4307_6740# 9.94e-21
C811 a_2376_6263# _03_ 0.171893f
C812 net11 a_4903_6575# 9.19e-19
C813 a_5547_7119# _02_ 0.001342f
C814 n_d[2] n_d[1] 0.157782f
C815 _09_ a_3057_6147# 2.03e-19
C816 net1 net7 0.002205f
C817 _09_ a_3111_5639# 0.101173f
C818 n_d[0] y_d[4] 0.002664f
C819 a_5476_6351# _02_ 4.67e-19
C820 a_4031_6740# a_4028_5467# 0.001113f
C821 net17 a_3859_7379# 0.006731f
C822 a_2376_6263# net3 0.279513f
C823 a_3111_5639# a_2939_6549# 1.29e-19
C824 a_2667_3463# a_2737_3561# 0.011552f
C825 a_2869_6147# _02_ 1.5e-20
C826 net18 net2 8.4e-20
C827 net1 _00_ 0.08935f
C828 net14 _00_ 0.013192f
C829 net8 net4 0.005588f
C830 a_2607_6147# net2 2.87e-19
C831 net18 y_d[7] 0.047502f
C832 a_4903_6575# net6 1.13e-19
C833 y_d[0] _02_ 1.15e-20
C834 net18 y_d[6] 0.026882f
C835 y_d[5] a_3384_5467# 1.67e-20
C836 net16 _03_ 5.56e-20
C837 a_3057_6147# a_2975_6147# 0.004937f
C838 a_3219_3463# VPWR 0.173446f
C839 a_3619_6147# a_3615_4943# 5.49e-22
C840 a_2975_6147# a_3111_5639# 3.1e-20
C841 a_4745_5533# a_4779_7379# 4.99e-21
C842 n_d[1] a_3384_5467# 5.48e-22
C843 a_3513_6147# _03_ 0.032416f
C844 net3 net16 0.006205f
C845 a_4031_6740# net19 0.027332f
C846 a_3513_6147# net3 0.062176f
C847 a_2821_3561# VPWR 0.015293f
C848 y_d[4] a_3384_5467# 1.21e-19
C849 n_d[0] net19 0.247879f
C850 net3 a_4745_5533# 0.006386f
C851 a_5297_6147# net19 0.001986f
C852 _02_ a_2667_5175# 0.212015f
C853 a_3707_3311# _06_ 6.02e-19
C854 _02_ a_2387_4373# 0.02199f
C855 net1 a_3061_3971# 0.087489f
C856 in[1] VPWR 0.143158f
C857 a_4249_6147# net1 0.055756f
C858 VPWR a_3309_5309# 8.53e-20
C859 a_3111_5639# a_3342_5493# 0.004898f
C860 _02_ a_2879_2223# 7.47e-19
C861 _00_ a_6112_6351# 3.96e-19
C862 a_3019_7338# a_4399_7338# 7.18e-21
C863 n_d[6] net19 2.97e-22
C864 a_5687_6740# VPWR 0.242732f
C865 _09_ a_4031_6740# 5.01e-19
C866 net12 _02_ 0.13023f
C867 a_3111_5639# a_3155_5056# 2.11e-19
C868 a_2939_6549# a_4031_6740# 1.14e-19
C869 a_2511_6147# _03_ 8.76e-19
C870 a_4167_3311# _02_ 0.231872f
C871 a_4355_6147# a_4509_6147# 0.008535f
C872 a_3289_3561# VPWR 0.008753f
C873 VPWR a_6651_7119# 0.453222f
C874 a_5297_6147# net10 0.137659f
C875 a_2387_7379# net3 2.53e-20
C876 _09_ n_d[0] 0.022414f
C877 net11 a_4031_6740# 4.9e-20
C878 net8 a_4307_6740# 5.07e-19
C879 net13 a_2961_3855# 4.54e-20
C880 a_2511_6147# net3 0.002388f
C881 a_2607_6147# a_2376_6263# 0.004999f
C882 a_3513_6147# a_3619_6147# 0.13675f
C883 n_d[0] a_2939_6549# 0.332224f
C884 _09_ n_d[2] 0.091851f
C885 y_d[5] _04_ 9.92e-19
C886 a_3384_5467# net19 1.9e-20
C887 n_d[2] a_2939_6549# 5.39e-20
C888 net2 a_3571_4074# 0.036667f
C889 a_4779_7379# net7 0.24588f
C890 n_d[6] net10 0.022509f
C891 a_3057_6147# net1 8.49e-19
C892 net11 a_5297_6147# 2.88e-21
C893 n_d[1] _04_ 0.003494f
C894 a_4355_6147# net2 0.121938f
C895 _03_ net7 3.33e-20
C896 a_5297_6147# a_5560_6351# 0.010598f
C897 a_4399_7338# a_3307_7379# 1.14e-19
C898 _02_ net4 2.07e-19
C899 _07_ net17 6.05e-20
C900 _00_ a_4779_7379# 2.99e-19
C901 net3 net7 0.014806f
C902 n_d[7] net9 0.073915f
C903 a_4031_6740# net6 0.108887f
C904 net11 n_d[6] 1.86e-19
C905 _00_ _03_ 1.9e-20
C906 net2 _02_ 0.215335f
C907 a_2387_5461# a_3111_5639# 3.54e-19
C908 in[0] _02_ 9.78e-20
C909 a_4028_5467# _04_ 1.42e-19
C910 net3 _00_ 0.534506f
C911 n_d[0] net6 4.66e-19
C912 a_5297_6147# _10_ 0.004189f
C913 a_3755_5639# net4 4.47e-22
C914 a_3384_5467# a_2939_6549# 9.7e-21
C915 a_2387_3027# a_2961_2767# 8.4e-20
C916 VPWR a_5849_6147# 0.147761f
C917 n_d[2] net6 0.024445f
C918 y_d[5] VPWR 0.559654f
C919 net8 a_4745_5533# 1.69e-20
C920 a_3129_6147# net2 1.42e-19
C921 net8 net9 0.007994f
C922 net2 a_3755_5639# 3.95e-19
C923 n_d[1] VPWR 0.966135f
C924 y_d[5] a_3491_6549# 0.328692f
C925 y_d[1] y_d[0] 0.091646f
C926 a_5547_7119# a_6099_7119# 0.003298f
C927 y_d[4] VPWR 0.514531f
C928 n_d[1] a_3491_6549# 1.62e-19
C929 a_2387_7379# net18 0.294339f
C930 net19 _04_ 0.021751f
C931 n_d[3] net7 0.02329f
C932 a_4355_6147# a_4307_6740# 1.4e-19
C933 a_4249_6147# _03_ 0.044411f
C934 _00_ a_2961_3855# 0.169071f
C935 a_3619_6147# _00_ 7.52e-22
C936 a_3219_3463# a_3289_3561# 0.011552f
C937 net3 a_3061_3971# 5.49e-21
C938 VPWR a_4028_5467# 0.203222f
C939 net1 a_4031_6740# 8.86e-20
C940 a_4249_6147# net3 0.095409f
C941 n_d[3] _00_ 3.78e-22
C942 _08_ a_3307_7379# 4.39e-20
C943 a_4443_3855# net1 3.31e-19
C944 a_4903_6575# a_4779_7379# 0.010769f
C945 _02_ a_3615_4943# 0.036642f
C946 n_d[7] net7 2.94e-20
C947 net1 _06_ 0.116701f
C948 n_d[0] net1 1.5e-19
C949 a_4903_6575# _03_ 1.97e-19
C950 a_5297_6147# net1 2.24e-19
C951 _02_ a_4307_6740# 1.45e-19
C952 VPWR a_2821_4943# 0.015734f
C953 _08_ a_3261_5493# 3.82e-19
C954 a_3384_5467# a_3342_5493# 1.84e-19
C955 a_4437_6147# _04_ 9.18e-19
C956 a_3755_5639# a_3905_5493# 0.002605f
C957 y_d[1] a_2879_2223# 7.91e-21
C958 _09_ _04_ 0.007929f
C959 VPWR a_2387_2197# 0.401728f
C960 a_2939_6549# _04_ 4.13e-19
C961 n_d[1] net5 0.027133f
C962 y_d[1] net12 0.003088f
C963 _08_ a_2667_5175# 3.66e-20
C964 a_3384_5467# a_3155_5056# 7.21e-19
C965 a_3755_5639# a_3615_4943# 0.01047f
C966 net4 _05_ 0.18294f
C967 n_d[0] a_2387_5461# 1.16e-21
C968 VPWR net19 0.285907f
C969 a_2387_3027# VPWR 0.438914f
C970 a_5547_7119# n_d[4] 0.356223f
C971 a_3111_5639# _03_ 3.35e-21
C972 net8 net7 0.087425f
C973 net11 _04_ 1.52e-20
C974 a_2961_3855# a_3061_3971# 0.167615f
C975 net2 a_4399_7338# 1.61e-20
C976 a_5353_6575# net19 7.47e-19
C977 a_3307_7379# a_3859_7379# 0.003298f
C978 a_3707_3311# VPWR 0.272595f
C979 a_3057_6147# net3 0.002054f
C980 a_3619_6147# a_4249_6147# 8.06e-19
C981 a_2387_3027# net15 1.19e-21
C982 net2 _05_ 0.029195f
C983 net3 a_3111_5639# 0.246257f
C984 a_3148_4215# net2 1.62e-20
C985 y_d[7] a_4399_7338# 1.44e-19
C986 a_3491_6549# net19 0.041342f
C987 a_2975_6147# _04_ 0.101833f
C988 net8 _00_ 0.047644f
C989 a_3701_6147# net1 8.93e-20
C990 a_5547_7119# n_d[5] 3.78e-19
C991 net1 a_3384_5467# 0.00111f
C992 net16 _02_ 0.096151f
C993 VPWR a_4437_6147# 1.73e-19
C994 a_3513_6147# _02_ 2.54e-21
C995 VPWR net10 0.816554f
C996 _04_ net6 0.025804f
C997 net13 _02_ 0.086326f
C998 _09_ VPWR 0.494198f
C999 a_4745_5533# _02_ 0.110884f
C1000 _02_ net9 0.001892f
C1001 n_d[3] a_4903_6575# 8.45e-20
C1002 VPWR a_2939_6549# 0.424108f
C1003 a_3773_6147# net17 8.47e-19
C1004 y_d[1] in[0] 0.320536f
C1005 y_d[0] y_d[2] 3.32e-20
C1006 net16 a_3755_5639# 1.75e-21
C1007 _09_ a_3491_6549# 0.007046f
C1008 net11 VPWR 1.00501f
C1009 a_2939_6549# a_3491_6549# 0.003298f
C1010 net11 a_5353_6575# 0.010835f
C1011 net19 net5 4.59e-20
C1012 _08_ net4 1.46e-20
C1013 VPWR a_5560_6351# 0.002658f
C1014 a_3155_5056# _04_ 4.51e-21
C1015 VPWR a_2975_6147# 0.128399f
C1016 a_4307_6740# a_4399_7338# 1.44e-19
C1017 net2 _08_ 0.036841f
C1018 _05_ a_4307_6740# 0.032822f
C1019 a_4031_6740# _03_ 0.00298f
C1020 a_4355_6147# net7 0.001361f
C1021 VPWR net6 0.54819f
C1022 a_2667_3463# a_2879_2223# 5.14e-20
C1023 VPWR _10_ 1.4496f
C1024 net3 a_4031_6740# 3.15e-19
C1025 net8 a_4903_6575# 0.115706f
C1026 n_d[0] _03_ 5.26e-21
C1027 n_d[2] a_4779_7379# 1.05e-21
C1028 a_4443_3855# net3 0.251966f
C1029 a_5297_6147# _03_ 1.16e-19
C1030 _09_ net5 4.42e-20
C1031 net1 _04_ 0.684292f
C1032 _00_ a_3571_4074# 0.002983f
C1033 a_2667_3463# net12 2.12e-21
C1034 a_4355_6147# _00_ 4.72e-21
C1035 y_d[2] net12 8.47e-19
C1036 net3 _06_ 0.002914f
C1037 net4 a_3859_7379# 1.43e-19
C1038 a_3491_6549# net6 0.234064f
C1039 _10_ a_3491_6549# 4.55e-20
C1040 n_d[0] net3 0.001282f
C1041 a_5297_6147# net3 8.24e-20
C1042 a_3219_3463# a_3707_3311# 0.117912f
C1043 n_d[2] net3 1.56e-21
C1044 _02_ net7 0.349514f
C1045 a_2667_5175# a_3237_5309# 3.04e-19
C1046 net2 a_3859_7379# 9.7e-20
C1047 net17 a_3261_5493# 1.08e-20
C1048 VPWR a_3155_5056# 0.181272f
C1049 _08_ a_3905_5493# 2.91e-20
C1050 _00_ _02_ 3.04333f
C1051 y_d[7] a_3859_7379# 2.94e-19
C1052 net15 a_3155_5056# 6.44e-20
C1053 VPWR a_3431_2223# 0.246601f
C1054 net17 a_2667_5175# 6.8e-21
C1055 a_3513_6147# _05_ 5.72e-19
C1056 _08_ a_3615_4943# 0.201372f
C1057 a_3148_4215# net13 3.22e-21
C1058 a_3384_5467# _03_ 3.72e-20
C1059 a_3061_3971# a_3571_4074# 0.01869f
C1060 a_2961_3855# _06_ 0.001326f
C1061 a_3129_6147# _00_ 1.75e-20
C1062 net6 net5 0.002356f
C1063 a_5687_6740# net19 0.108611f
C1064 _00_ a_3755_5639# 3.79e-19
C1065 net1 VPWR 3.48707f
C1066 net14 VPWR 0.401235f
C1067 a_4249_6147# a_4355_6147# 0.13675f
C1068 a_3701_6147# net3 0.002474f
C1069 net3 a_3384_5467# 0.063454f
C1070 n_d[1] y_d[5] 0.006272f
C1071 net14 net15 6.68e-20
C1072 a_2667_3463# in[0] 4.36e-21
C1073 y_d[2] in[0] 0.024732f
C1074 net1 net15 0.030091f
C1075 net1 a_3491_6549# 0.011058f
C1076 a_3289_3561# a_3707_3311# 2.64e-19
C1077 n_d[2] n_d[3] 0.084983f
C1078 y_d[5] y_d[4] 0.093893f
C1079 _02_ a_3061_3971# 0.002683f
C1080 VPWR a_2387_5461# 0.482421f
C1081 a_4249_6147# _02_ 3.76e-19
C1082 y_d[1] net13 0.026346f
C1083 a_5687_6740# net10 0.035637f
C1084 a_2387_5461# net15 2.69e-21
C1085 net10 a_6651_7119# 1.79e-19
C1086 net16 _08_ 9.79e-20
C1087 a_7111_6575# net9 0.011283f
C1088 net2 a_3237_5309# 4.89e-19
C1089 n_d[1] a_4028_5467# 1.35e-20
C1090 net18 n_d[2] 0.014524f
C1091 n_d[7] n_d[6] 0.113801f
C1092 net4 net17 0.042705f
C1093 a_3701_6147# a_3619_6147# 0.004937f
C1094 a_3513_6147# _08_ 9.44e-19
C1095 net11 a_5687_6740# 0.024027f
C1096 a_4903_6575# _02_ 0.014136f
C1097 y_d[4] a_4028_5467# 2.01e-20
C1098 VPWR a_6112_6351# 0.001755f
C1099 _04_ a_4779_7379# 0.021795f
C1100 net1 net5 1.5e-21
C1101 a_4399_7338# net7 7.82e-20
C1102 net8 a_5297_6147# 3.06e-19
C1103 net2 net17 0.045229f
C1104 a_6099_7119# net9 0.028688f
C1105 _03_ _04_ 0.222355f
C1106 net11 a_6651_7119# 0.002354f
C1107 _07_ net4 1.76e-19
C1108 y_d[7] net17 2.43e-36
C1109 y_d[5] net19 0.32326f
C1110 a_3111_5639# _02_ 0.001539f
C1111 net3 _04_ 0.41588f
C1112 net8 n_d[6] 6.07e-20
C1113 a_3148_4215# _00_ 3.71e-20
C1114 n_d[1] net19 7.59e-21
C1115 in[2] VPWR 0.264075f
C1116 net2 _07_ 0.001497f
C1117 y_d[0] a_3045_2767# 6.6e-21
C1118 a_5687_6740# _10_ 0.189829f
C1119 VPWR a_3986_5493# 4.09e-20
C1120 a_3219_3463# net1 0.012321f
C1121 a_3111_5639# a_3755_5639# 1.56e-19
C1122 a_5849_6147# net10 0.126485f
C1123 a_2667_5175# a_2737_4943# 0.011552f
C1124 a_3155_5056# a_3309_5309# 0.004009f
C1125 _09_ y_d[5] 0.035382f
C1126 VPWR a_4779_7379# 0.461185f
C1127 a_4028_5467# net19 1.7e-20
C1128 in[1] a_3431_2223# 7.6e-20
C1129 y_d[5] a_2939_6549# 0.152546f
C1130 _09_ n_d[1] 0.071967f
C1131 VPWR _03_ 0.422323f
C1132 net14 a_2821_3561# 0.002266f
C1133 a_3619_6147# _04_ 0.041068f
C1134 n_d[4] net9 9.12e-20
C1135 n_d[1] a_2939_6549# 2.16e-19
C1136 net17 a_3615_4943# 0.109442f
C1137 net11 a_5849_6147# 0.001219f
C1138 net3 VPWR 2.68627f
C1139 n_d[3] _04_ 0.026471f
C1140 a_4249_6147# _05_ 0.007929f
C1141 _09_ y_d[4] 0.001269f
C1142 a_3148_4215# a_3061_3971# 0.004898f
C1143 net17 a_4307_6740# 4.59e-19
C1144 a_3019_7338# a_3307_7379# 0.001856f
C1145 a_3491_6549# _03_ 2.62e-19
C1146 in[1] net1 1.61e-19
C1147 a_2667_3463# net13 0.119585f
C1148 a_3571_4074# _06_ 0.216565f
C1149 net3 net15 9.12e-20
C1150 y_d[2] net13 3.96e-20
C1151 net12 a_3045_2767# 0.016223f
C1152 a_2387_3027# a_2387_2197# 0.050529f
C1153 net3 a_3491_6549# 3.95e-19
C1154 _00_ _08_ 0.09833f
C1155 n_d[5] net9 0.026309f
C1156 _02_ a_4031_6740# 7.96e-20
C1157 _07_ a_4307_6740# 2.37e-19
C1158 net13 a_2737_3561# 2.64e-19
C1159 a_3289_3561# net1 0.001023f
C1160 net16 a_3237_5309# 2.01e-20
C1161 y_d[5] net6 0.035657f
C1162 a_5849_6147# _10_ 0.020602f
C1163 _02_ _06_ 3.08e-19
C1164 a_5297_6147# _02_ 0.155083f
C1165 n_d[1] net6 0.084018f
C1166 a_4779_7379# net5 0.001473f
C1167 VPWR a_2961_3855# 0.193136f
C1168 a_3619_6147# VPWR 0.130415f
C1169 _03_ net5 4.75e-21
C1170 net16 net17 5.05e-19
C1171 a_3755_5639# a_4031_6740# 1.54e-20
C1172 net8 _04_ 0.001321f
C1173 n_d[3] VPWR 0.460331f
C1174 net15 a_2961_3855# 0.002394f
C1175 net10 net19 0.010531f
C1176 _09_ net19 0.03154f
C1177 net3 net5 9.7e-19
C1178 a_3513_6147# net17 0.005185f
C1179 a_3619_6147# a_3491_6549# 0.001225f
C1180 a_2939_6549# net19 0.056677f
C1181 y_d[3] VPWR 0.505033f
C1182 net4 a_2387_6549# 3.32e-19
C1183 a_2869_6147# a_2667_5175# 4.74e-20
C1184 a_4028_5467# net6 9.92e-22
C1185 n_d[4] net7 0.002262f
C1186 y_d[4] a_3342_5493# 3.47e-20
C1187 n_d[7] VPWR 0.628106f
C1188 y_d[3] net15 0.02628f
C1189 net11 net19 0.207115f
C1190 net2 a_2387_6549# 0.011173f
C1191 n_d[4] _00_ 8.69e-19
C1192 net18 VPWR 0.195526f
C1193 a_4745_5533# _07_ 3.43e-19
C1194 _10_ a_5008_5487# 3.89e-19
C1195 a_3384_5467# _02_ 0.003683f
C1196 y_d[7] a_2387_6549# 0.397458f
C1197 _10_ a_2821_4943# 2.49e-20
C1198 a_2975_6147# net19 1.68e-20
C1199 a_2607_6147# VPWR 0.001803f
C1200 net1 a_5849_6147# 3.43e-20
C1201 y_d[5] net1 1.88e-19
C1202 a_2667_3463# _00_ 0.072341f
C1203 y_d[0] a_2879_2223# 0.337682f
C1204 y_d[6] a_2387_6549# 8.94e-19
C1205 _09_ a_2939_6549# 0.038262f
C1206 n_d[1] net1 5.45e-19
C1207 net8 VPWR 0.668331f
C1208 a_3773_6147# net2 9.85e-19
C1209 net11 net10 0.043875f
C1210 net8 a_5353_6575# 5.2e-19
C1211 net19 net6 0.016964f
C1212 _10_ net19 0.00313f
C1213 y_d[0] net12 0.049027f
C1214 n_d[3] net5 0.008654f
C1215 a_3111_5639# _08_ 0.002261f
C1216 a_3755_5639# a_3384_5467# 9.28e-19
C1217 y_d[4] net1 7.19e-19
C1218 a_5560_6351# net10 0.005356f
C1219 a_2667_5175# a_2387_4373# 6.46e-19
C1220 a_3019_7338# y_d[7] 0.010978f
C1221 _09_ a_2975_6147# 0.013436f
C1222 a_4031_6740# _05_ 0.213819f
C1223 _00_ a_3237_5309# 8.4e-19
C1224 _02_ a_2961_2767# 9.04e-19
C1225 net1 a_4028_5467# 0.081631f
C1226 a_2975_6147# a_2939_6549# 0.001159f
C1227 a_3019_7338# y_d[6] 9.24e-20
C1228 a_4355_6147# _04_ 0.048879f
C1229 net17 net7 1.34e-20
C1230 y_d[4] a_2387_5461# 0.341222f
C1231 _00_ a_5437_6575# 1.5e-19
C1232 n_d[0] _05_ 8.92e-21
C1233 n_d[2] a_4399_7338# 1.18e-19
C1234 _10_ net10 0.228061f
C1235 net18 net5 0.002326f
C1236 _09_ net6 0.054062f
C1237 net2 a_2869_6147# 0.135865f
C1238 net12 a_2879_2223# 0.23376f
C1239 net4 a_3307_7379# 0.00683f
C1240 a_2939_6549# net6 0.002256f
C1241 _00_ net17 0.020938f
C1242 a_5849_6147# a_6112_6351# 0.010598f
C1243 net14 a_2387_2197# 1.11e-19
C1244 y_d[7] a_2869_6147# 4.79e-20
C1245 net1 a_2387_2197# 2.53e-19
C1246 a_2376_6263# a_2387_6549# 0.011645f
C1247 _07_ net7 0.039702f
C1248 _02_ _04_ 3.64e-19
C1249 net11 net6 0.001335f
C1250 net2 a_3307_7379# 0.001163f
C1251 net11 _10_ 0.004176f
C1252 net8 net5 7.76e-21
C1253 y_d[0] net2 9.23e-20
C1254 y_d[0] in[0] 0.201175f
C1255 a_2387_3027# net14 0.2058f
C1256 net1 net19 6.53e-19
C1257 net16 a_2737_4943# 0.00346f
C1258 _00_ _07_ 0.009575f
C1259 _09_ a_3155_5056# 3.85e-19
C1260 a_3707_3311# net1 0.23412f
C1261 y_d[7] a_3307_7379# 9.06e-19
C1262 net2 a_3261_5493# 8.89e-19
C1263 a_3129_6147# _04_ 7.69e-20
C1264 a_2939_6549# a_3155_5056# 2.15e-21
C1265 VPWR a_3571_4074# 0.2678f
C1266 a_4745_5533# a_4924_5487# 0.007688f
C1267 a_4355_6147# VPWR 0.150289f
C1268 net16 a_2387_6549# 4.71e-21
C1269 net15 a_3571_4074# 0.108671f
C1270 a_2387_5461# net19 2.08e-20
C1271 net13 a_3045_2767# 4.85e-19
C1272 net2 a_2667_5175# 0.005158f
C1273 net2 a_2387_4373# 2.98e-19
C1274 net1 net10 9.89e-21
C1275 net1 a_4437_6147# 0.002177f
C1276 a_4249_6147# net17 5.08e-19
C1277 _08_ _06_ 8.23e-20
C1278 net13 a_3373_3561# 0.002266f
C1279 net2 a_2879_2223# 1.4e-19
C1280 _09_ net1 0.025471f
C1281 in[0] a_2879_2223# 0.104281f
C1282 a_2975_6147# a_3155_5056# 2.02e-21
C1283 VPWR _02_ 2.19337f
C1284 n_d[6] a_7111_6575# 0.345034f
C1285 net1 a_2939_6549# 6.05e-20
C1286 y_d[4] a_3986_5493# 3.68e-21
C1287 n_d[1] a_4779_7379# 1.98e-19
C1288 a_5353_6575# _02_ 5.37e-19
C1289 net12 net2 9.15e-21
C1290 y_d[5] net3 5.52e-19
C1291 in[0] net12 0.126451f
C1292 _02_ net15 0.030359f
C1293 a_4249_6147# _07_ 5.72e-19
C1294 a_4167_3311# net2 0.245173f
C1295 _02_ a_3491_6549# 2.3e-20
C1296 a_2376_6263# a_2869_6147# 0.001158f
C1297 a_4903_6575# net17 9.72e-20
C1298 _10_ a_3155_5056# 0.092458f
C1299 _09_ a_2387_5461# 0.048064f
C1300 a_4028_5467# a_3986_5493# 1.84e-19
C1301 n_d[1] net3 5.57e-20
C1302 n_d[7] a_6651_7119# 0.145199f
C1303 y_d[4] _03_ 0.002691f
C1304 a_4031_6740# a_3859_7379# 0.011387f
C1305 a_6099_7119# n_d[6] 2.2e-19
C1306 a_3129_6147# VPWR 1.64e-19
C1307 VPWR a_3755_5639# 0.203377f
C1308 net1 a_2975_6147# 0.048721f
C1309 y_d[4] net3 9.5e-19
C1310 a_2387_7379# a_2387_6549# 0.050529f
C1311 _07_ a_4903_6575# 0.193402f
C1312 _03_ a_4028_5467# 6.96e-20
C1313 a_4509_6147# net2 2.44e-19
C1314 net8 a_5687_6740# 0.046967f
C1315 a_3755_5639# a_3491_6549# 1.55e-21
C1316 a_3111_5639# net17 5.31e-20
C1317 a_3701_6147# _08_ 1.18e-19
C1318 a_3384_5467# _08_ 0.012436f
C1319 n_d[2] a_3859_7379# 8.25e-19
C1320 a_4399_7338# _04_ 0.197382f
C1321 net1 net6 9.97e-20
C1322 a_4924_5487# net7 0.001923f
C1323 a_6112_6351# net10 7.31e-19
C1324 net1 _10_ 0.020959f
C1325 net2 net4 7.75e-19
C1326 net3 a_4028_5467# 0.028208f
C1327 _05_ _04_ 0.023652f
C1328 _02_ net5 6.22e-20
C1329 _00_ a_4924_5487# 0.001001f
C1330 y_d[7] net4 0.003786f
C1331 a_2376_6263# a_2667_5175# 4.55e-20
C1332 net3 a_5008_5487# 5.52e-19
C1333 n_d[4] a_5297_6147# 1.32e-21
C1334 n_d[1] a_3619_6147# 6.31e-20
C1335 in[0] net2 5.95e-22
C1336 a_2387_7379# a_3019_7338# 0.001557f
C1337 net19 a_4779_7379# 1.3e-19
C1338 net11 a_6112_6351# 5.87e-20
C1339 _00_ a_3045_2767# 3.34e-19
C1340 y_d[7] net2 0.005273f
C1341 a_3219_3463# a_3571_4074# 3.14e-19
C1342 n_d[1] n_d[3] 0.001222f
C1343 net1 a_3155_5056# 0.002438f
C1344 _03_ net19 0.048018f
C1345 a_3373_3561# _00_ 0.002384f
C1346 n_d[4] n_d[6] 7.01e-20
C1347 y_d[0] net13 0.08809f
C1348 net3 net19 0.001032f
C1349 net1 a_3431_2223# 0.110108f
C1350 y_d[6] y_d[7] 0.073731f
C1351 y_d[4] y_d[3] 0.092925f
C1352 VPWR a_4399_7338# 0.267703f
C1353 net16 a_2667_5175# 0.150346f
C1354 a_3219_3463# _02_ 0.185099f
C1355 net16 a_2387_4373# 0.002198f
C1356 net18 n_d[1] 0.132961f
C1357 n_d[5] n_d[6] 0.162825f
C1358 a_6112_6351# _10_ 0.001393f
C1359 VPWR _05_ 0.260037f
C1360 net14 net1 8.54e-20
C1361 a_3148_4215# VPWR 4.38e-20
C1362 a_4437_6147# _03_ 2.83e-19
C1363 y_d[0] VGND 2.03303f
C1364 y_d[1] VGND 1.1568f
C1365 in[2] VGND 1.55542f
C1366 in[1] VGND 1.44541f
C1367 in[0] VGND 1.29688f
C1368 y_d[2] VGND 1.214f
C1369 y_d[3] VGND 1.24123f
C1370 y_d[4] VGND 1.22235f
C1371 n_d[6] VGND 1.39038f
C1372 y_d[5] VGND 0.986898f
C1373 n_d[0] VGND 2.40927f
C1374 y_d[7] VGND 1.82189f
C1375 n_d[5] VGND 1.09526f
C1376 n_d[7] VGND 2.46115f
C1377 n_d[4] VGND 1.17565f
C1378 n_d[3] VGND 1.30988f
C1379 n_d[1] VGND 1.25545f
C1380 n_d[2] VGND 1.12337f
C1381 y_d[6] VGND 1.22055f
C1382 VPWR VGND 0.151325p
C1383 a_7437_2388# VGND 0.292925f
C1384 a_5137_2388# VGND 0.29556f
C1385 a_3431_2223# VGND 0.31543f
C1386 a_2879_2223# VGND 0.561941f
C1387 a_2387_2197# VGND 0.560962f
C1388 a_3045_2767# VGND 4.15e-19
C1389 a_2961_2767# VGND 3.93e-19
C1390 net12 VGND 0.367348f
C1391 a_2387_3027# VGND 0.555755f
C1392 a_3373_3561# VGND 0.005743f
C1393 a_3289_3561# VGND 0.001255f
C1394 net13 VGND 0.835782f
C1395 a_2821_3561# VGND 5.29e-19
C1396 a_2737_3561# VGND 8.02e-19
C1397 net14 VGND 0.695731f
C1398 a_4167_3311# VGND 0.333021f
C1399 a_3707_3311# VGND 0.330291f
C1400 a_3219_3463# VGND 0.22679f
C1401 a_2667_3463# VGND 0.222207f
C1402 a_3220_4215# VGND 0.00266f
C1403 a_3148_4215# VGND 4.66e-19
C1404 a_4443_3855# VGND 0.353009f
C1405 _06_ VGND 0.302728f
C1406 a_3571_4074# VGND 0.272309f
C1407 a_3061_3971# VGND 0.245958f
C1408 a_2961_3855# VGND 0.211241f
C1409 net15 VGND 0.846618f
C1410 a_2387_4373# VGND 0.62901f
C1411 a_2821_4943# VGND 7.16e-20
C1412 a_2737_4943# VGND 8.99e-19
C1413 a_3309_5309# VGND 0.002704f
C1414 a_3237_5309# VGND 7.03e-19
C1415 a_3615_4943# VGND 0.251104f
C1416 a_3155_5056# VGND 0.273669f
C1417 a_2667_5175# VGND 0.207107f
C1418 a_5008_5487# VGND 0.012872f
C1419 a_4924_5487# VGND 0.009823f
C1420 a_3986_5493# VGND 4.85e-19
C1421 a_3905_5493# VGND 0.002577f
C1422 a_3342_5493# VGND 0.001171f
C1423 a_3261_5493# VGND 0.003377f
C1424 a_4028_5467# VGND 0.202544f
C1425 a_4745_5533# VGND 0.325283f
C1426 _08_ VGND 0.460475f
C1427 a_3384_5467# VGND 0.240632f
C1428 a_3755_5639# VGND 0.226791f
C1429 a_3111_5639# VGND 0.276648f
C1430 net16 VGND 0.728393f
C1431 a_2387_5461# VGND 0.561079f
C1432 a_4509_6147# VGND 1.72e-19
C1433 a_4437_6147# VGND 1.19e-19
C1434 a_3773_6147# VGND 2.07e-19
C1435 a_3701_6147# VGND 1.32e-19
C1436 a_3129_6147# VGND 1.25e-19
C1437 a_3057_6147# VGND 8.48e-20
C1438 a_6112_6351# VGND 0.009062f
C1439 a_6028_6351# VGND 0.006966f
C1440 a_5560_6351# VGND 0.006912f
C1441 a_5476_6351# VGND 0.005722f
C1442 a_5849_6147# VGND 0.287754f
C1443 a_5297_6147# VGND 0.296838f
C1444 a_4355_6147# VGND 0.365445f
C1445 a_4249_6147# VGND 0.218144f
C1446 a_3619_6147# VGND 0.351049f
C1447 a_3513_6147# VGND 0.227181f
C1448 a_2975_6147# VGND 0.330936f
C1449 a_2869_6147# VGND 0.207257f
C1450 net2 VGND 2.70606f
C1451 net1 VGND 1.6913f
C1452 net3 VGND 4.42304f
C1453 a_2376_6263# VGND 0.359054f
C1454 a_5437_6575# VGND 5.32e-19
C1455 a_5353_6575# VGND 5.3e-19
C1456 a_7111_6575# VGND 0.62073f
C1457 net10 VGND 1.12948f
C1458 _10_ VGND 1.20229f
C1459 a_5687_6740# VGND 0.263586f
C1460 _00_ VGND 3.19786f
C1461 _02_ VGND 3.41078f
C1462 a_4903_6575# VGND 0.270408f
C1463 _07_ VGND 0.512249f
C1464 _03_ VGND 0.962736f
C1465 a_4307_6740# VGND 0.233816f
C1466 _05_ VGND 0.353103f
C1467 a_4031_6740# VGND 0.206347f
C1468 net17 VGND 0.554795f
C1469 a_3491_6549# VGND 0.548212f
C1470 net4 VGND 0.264102f
C1471 a_2939_6549# VGND 0.563756f
C1472 net19 VGND 1.77539f
C1473 a_2387_6549# VGND 0.54012f
C1474 a_6651_7119# VGND 0.624828f
C1475 net9 VGND 1.16017f
C1476 a_6099_7119# VGND 0.69196f
C1477 net11 VGND 0.475474f
C1478 a_5547_7119# VGND 0.605951f
C1479 net8 VGND 0.409176f
C1480 net7 VGND 0.655417f
C1481 a_4779_7379# VGND 0.719039f
C1482 _04_ VGND 0.418939f
C1483 a_4399_7338# VGND 0.261742f
C1484 net5 VGND 0.36733f
C1485 a_3859_7379# VGND 0.559281f
C1486 net6 VGND 0.325689f
C1487 a_3307_7379# VGND 0.628211f
C1488 _09_ VGND 0.459189f
C1489 a_3019_7338# VGND 0.242623f
C1490 net18 VGND 0.376089f
C1491 a_2387_7379# VGND 0.56939f
C1492 _01_.n0 VGND 0.675402f
C1493 _01_.t0 VGND 0.029635f
C1494 _01_.t1 VGND 0.029635f
C1495 _01_.n1 VGND 0.061446f
C1496 _01_.t12 VGND 0.049941f
C1497 _01_.t20 VGND 0.03136f
C1498 _01_.n2 VGND 0.067522f
C1499 _37_.B VGND 0.124687f
C1500 _01_.t11 VGND 0.020075f
C1501 _01_.t5 VGND 0.021519f
C1502 _01_.n3 VGND 0.062647f
C1503 _34_.A_N VGND 0.045419f
C1504 _01_.t14 VGND 0.031029f
C1505 _01_.t21 VGND 0.049535f
C1506 _01_.n4 VGND 0.076763f
C1507 _31_.B VGND 0.013401f
C1508 _01_.n5 VGND 0.080296f
C1509 _25_.B VGND 0.019197f
C1510 _01_.t16 VGND 0.049535f
C1511 _01_.t6 VGND 0.031029f
C1512 _01_.n6 VGND 0.076564f
C1513 _01_.n7 VGND 0.041034f
C1514 _01_.n8 VGND 0.333909f
C1515 _32_.A_N VGND 0.084586f
C1516 _01_.t7 VGND 0.027479f
C1517 _01_.t19 VGND 0.019773f
C1518 _01_.n9 VGND 0.025376f
C1519 _01_.n10 VGND 0.0734f
C1520 _01_.n11 VGND 0.082816f
C1521 _01_.n12 VGND 0.025376f
C1522 _01_.n13 VGND 0.460769f
C1523 _01_.t9 VGND 0.03136f
C1524 _01_.t15 VGND 0.049941f
C1525 _01_.n14 VGND 0.068055f
C1526 _26_.A VGND 0.124762f
C1527 _01_.t4 VGND 0.047328f
C1528 _01_.t18 VGND 0.08663f
C1529 _35_.B VGND 0.08726f
C1530 _01_.n15 VGND 0.445407f
C1531 _01_.n16 VGND 0.484584f
C1532 _01_.t23 VGND 0.026892f
C1533 _01_.t22 VGND 0.020329f
C1534 _01_.n17 VGND 0.0591f
C1535 _17_.C_N VGND 0.011568f
C1536 _01_.n18 VGND 0.153387f
C1537 _01_.n19 VGND 0.412712f
C1538 _20_.B VGND 0.014488f
C1539 _01_.t8 VGND 0.049941f
C1540 _01_.t13 VGND 0.03136f
C1541 _01_.n20 VGND 0.067135f
C1542 _01_.n21 VGND 0.031503f
C1543 _01_.t10 VGND 0.03136f
C1544 _01_.t17 VGND 0.049941f
C1545 _01_.n22 VGND 0.074476f
C1546 _14_.B VGND 0.186381f
C1547 _01_.n23 VGND 0.541568f
C1548 _01_.n24 VGND 0.218907f
C1549 _01_.n25 VGND 0.085915f
C1550 _01_.t2 VGND 0.012446f
C1551 _01_.t3 VGND 0.012446f
C1552 _01_.n26 VGND 0.030677f
C1553 _12_.X VGND 0.230985f
C1554 VPWR.n0 VGND 0.001122f
C1555 VPWR.n1 VGND 8.79e-19
C1556 VPWR.n2 VGND 0.001099f
C1557 VPWR.n3 VGND 0.00196f
C1558 VPWR.n4 VGND 0.206033f
C1559 VPWR.n5 VGND 5.17e-19
C1560 VPWR.t93 VGND 0.004392f
C1561 VPWR.n6 VGND 0.005263f
C1562 VPWR.t87 VGND 0.001039f
C1563 VPWR.t89 VGND 0.001039f
C1564 VPWR.n7 VGND 0.002108f
C1565 VPWR.n8 VGND 0.001846f
C1566 VPWR.n9 VGND 0.003278f
C1567 VPWR.t252 VGND 0.003052f
C1568 VPWR.n10 VGND 0.002326f
C1569 VPWR.t91 VGND 0.00141f
C1570 VPWR.t360 VGND 0.001039f
C1571 VPWR.n11 VGND 0.002603f
C1572 VPWR.t533 VGND 0.040428f
C1573 VPWR.n12 VGND 0.018883f
C1574 VPWR.n13 VGND 0.003278f
C1575 VPWR.t321 VGND 0.004348f
C1576 VPWR.t315 VGND 0.001039f
C1577 VPWR.t317 VGND 0.001039f
C1578 VPWR.n14 VGND 0.002108f
C1579 VPWR.n15 VGND 0.003777f
C1580 VPWR.n16 VGND 0.003278f
C1581 VPWR.t319 VGND 0.00141f
C1582 VPWR.t59 VGND 0.001039f
C1583 VPWR.n17 VGND 0.002603f
C1584 VPWR.n18 VGND 0.002313f
C1585 VPWR.t467 VGND 0.004348f
C1586 VPWR.n19 VGND 0.005716f
C1587 VPWR.t253 VGND 0.003052f
C1588 VPWR.n20 VGND 0.002124f
C1589 VPWR.t278 VGND 8.5e-19
C1590 VPWR.t428 VGND 8.5e-19
C1591 VPWR.n21 VGND 0.001889f
C1592 VPWR.n22 VGND 0.004708f
C1593 VPWR.t469 VGND 0.001039f
C1594 VPWR.t463 VGND 0.001039f
C1595 VPWR.n23 VGND 0.002121f
C1596 VPWR.n24 VGND 0.001099f
C1597 VPWR.n25 VGND 0.00196f
C1598 VPWR.n26 VGND 0.263078f
C1599 VPWR.n27 VGND 0.001895f
C1600 VPWR.n28 VGND 0.001895f
C1601 VPWR.n29 VGND 0.129213f
C1602 VPWR.n30 VGND 0.00196f
C1603 VPWR.n31 VGND 3.05e-19
C1604 VPWR.n32 VGND 8.79e-19
C1605 VPWR.n33 VGND 0.001639f
C1606 VPWR.n34 VGND 0.004131f
C1607 VPWR.t39 VGND 0.00141f
C1608 VPWR.t388 VGND 0.001447f
C1609 VPWR.n35 VGND 0.00301f
C1610 VPWR.n36 VGND 0.005297f
C1611 VPWR.n37 VGND 0.003278f
C1612 VPWR.t55 VGND 6.35e-19
C1613 VPWR.t485 VGND 0.001025f
C1614 VPWR.n38 VGND 0.003075f
C1615 VPWR.t193 VGND 0.003052f
C1616 VPWR.n39 VGND 0.002371f
C1617 VPWR.n40 VGND 0.003288f
C1618 VPWR.n41 VGND 0.003278f
C1619 VPWR.t53 VGND 0.00141f
C1620 VPWR.t441 VGND 0.001447f
C1621 VPWR.n42 VGND 0.00301f
C1622 VPWR.t512 VGND 0.011578f
C1623 VPWR.t180 VGND 0.002774f
C1624 VPWR.n43 VGND 0.002735f
C1625 VPWR.n44 VGND 0.008976f
C1626 VPWR.n45 VGND 0.005383f
C1627 VPWR.t475 VGND 6.35e-19
C1628 VPWR.t392 VGND 0.001025f
C1629 VPWR.n46 VGND 0.003075f
C1630 VPWR.n47 VGND 0.00108f
C1631 VPWR.t128 VGND 0.036235f
C1632 VPWR.t443 VGND 0.025312f
C1633 VPWR.t415 VGND 0.009558f
C1634 VPWR.t413 VGND 0.009768f
C1635 VPWR.t24 VGND 0.009033f
C1636 VPWR.t419 VGND 0.010083f
C1637 VPWR.t365 VGND 0.009033f
C1638 VPWR.t417 VGND 0.007562f
C1639 VPWR.t13 VGND 0.003886f
C1640 VPWR.t353 VGND 0.009558f
C1641 VPWR.t366 VGND 0.009558f
C1642 VPWR.t429 VGND 0.024577f
C1643 VPWR.t16 VGND 0.009243f
C1644 VPWR.t421 VGND 0.009978f
C1645 VPWR.t28 VGND 0.009978f
C1646 VPWR.t34 VGND 0.010293f
C1647 VPWR.t425 VGND 0.009978f
C1648 VPWR.t21 VGND 0.010188f
C1649 VPWR.t267 VGND 0.011868f
C1650 VPWR.t19 VGND 0.01607f
C1651 VPWR.t301 VGND 0.012394f
C1652 VPWR.t439 VGND 0.014914f
C1653 VPWR.t362 VGND 0.009243f
C1654 VPWR.t96 VGND 0.009978f
C1655 VPWR.t26 VGND 0.009978f
C1656 VPWR.t30 VGND 0.010293f
C1657 VPWR.t451 VGND 0.009978f
C1658 VPWR.t363 VGND 0.010188f
C1659 VPWR.t289 VGND 0.012078f
C1660 VPWR.t389 VGND 0.006827f
C1661 VPWR.t32 VGND 0.003151f
C1662 VPWR.t490 VGND 0.011448f
C1663 VPWR.t116 VGND 0.007562f
C1664 VPWR.t23 VGND 0.013339f
C1665 VPWR.t372 VGND 0.015965f
C1666 VPWR.n48 VGND 0.012003f
C1667 VPWR.t373 VGND 6.39e-19
C1668 VPWR.t331 VGND 0.001002f
C1669 VPWR.n49 VGND 0.002906f
C1670 VPWR.t117 VGND 0.002797f
C1671 VPWR.n50 VGND 0.001637f
C1672 VPWR.n51 VGND 0.001817f
C1673 VPWR.t525 VGND 0.00583f
C1674 VPWR.n52 VGND 0.008822f
C1675 VPWR.n53 VGND 6.41e-19
C1676 VPWR.t390 VGND 0.001554f
C1677 VPWR.t33 VGND 0.001712f
C1678 VPWR.n54 VGND 0.001122f
C1679 VPWR.t290 VGND 4.21e-19
C1680 VPWR.t364 VGND 4.21e-19
C1681 VPWR.n55 VGND 8.5e-19
C1682 VPWR.n56 VGND 0.002972f
C1683 VPWR.n57 VGND 8.22e-19
C1684 VPWR.n58 VGND 0.003278f
C1685 VPWR.t27 VGND 6.39e-19
C1686 VPWR.t452 VGND 0.001002f
C1687 VPWR.n59 VGND 0.002948f
C1688 VPWR.n60 VGND 0.003278f
C1689 VPWR.t31 VGND 6.24e-19
C1690 VPWR.t97 VGND 2.58e-19
C1691 VPWR.n61 VGND 0.003251f
C1692 VPWR.t302 VGND 0.001554f
C1693 VPWR.n62 VGND 0.003525f
C1694 VPWR.n63 VGND 0.001942f
C1695 VPWR.t20 VGND 0.001698f
C1696 VPWR.n64 VGND 0.002458f
C1697 VPWR.t268 VGND 4.21e-19
C1698 VPWR.t22 VGND 4.21e-19
C1699 VPWR.n65 VGND 9.17e-19
C1700 VPWR.t29 VGND 6.39e-19
C1701 VPWR.t426 VGND 0.001002f
C1702 VPWR.n66 VGND 0.002948f
C1703 VPWR.n67 VGND 0.003278f
C1704 VPWR.n68 VGND 0.003278f
C1705 VPWR.t35 VGND 6.24e-19
C1706 VPWR.t422 VGND 2.58e-19
C1707 VPWR.n69 VGND 0.003251f
C1708 VPWR.n70 VGND 0.001161f
C1709 VPWR.n71 VGND 4.48e-19
C1710 VPWR.t367 VGND 0.001712f
C1711 VPWR.n72 VGND 6.24e-19
C1712 VPWR.n73 VGND 0.001104f
C1713 VPWR.t354 VGND 0.001039f
C1714 VPWR.t418 VGND 0.00141f
C1715 VPWR.n74 VGND 0.002645f
C1716 VPWR.t420 VGND 0.001039f
C1717 VPWR.t414 VGND 0.001039f
C1718 VPWR.n75 VGND 0.002121f
C1719 VPWR.n76 VGND 0.002973f
C1720 VPWR.n77 VGND 0.001176f
C1721 VPWR.n78 VGND 0.001099f
C1722 VPWR.n79 VGND 0.00196f
C1723 VPWR.n80 VGND 0.206033f
C1724 VPWR.n81 VGND 0.001895f
C1725 VPWR.n82 VGND 0.129213f
C1726 VPWR.n83 VGND 0.00196f
C1727 VPWR.n84 VGND 3.05e-19
C1728 VPWR.n85 VGND 8.79e-19
C1729 VPWR.t224 VGND 0.003052f
C1730 VPWR.n86 VGND 0.001069f
C1731 VPWR.n87 VGND 0.002458f
C1732 VPWR.t448 VGND 4.21e-19
C1733 VPWR.t473 VGND 4.21e-19
C1734 VPWR.n88 VGND 9.53e-19
C1735 VPWR.n89 VGND 0.00912f
C1736 VPWR.n90 VGND 0.003278f
C1737 VPWR.t397 VGND 6.24e-19
C1738 VPWR.t12 VGND -6.55e-19
C1739 VPWR.n91 VGND 0.004151f
C1740 VPWR.n92 VGND 0.004233f
C1741 VPWR.t546 VGND 0.040428f
C1742 VPWR.t57 VGND 8.5e-19
C1743 VPWR.t63 VGND 8.5e-19
C1744 VPWR.n93 VGND 0.001849f
C1745 VPWR.n94 VGND 0.007706f
C1746 VPWR.t159 VGND 0.003064f
C1747 VPWR.n95 VGND 0.00342f
C1748 VPWR.n96 VGND 0.001817f
C1749 VPWR.n97 VGND 0.011575f
C1750 VPWR.n98 VGND 0.001639f
C1751 VPWR.n99 VGND 0.001321f
C1752 VPWR.n100 VGND 8.79e-19
C1753 VPWR.n101 VGND 0.00196f
C1754 VPWR.n102 VGND 0.263078f
C1755 VPWR.n103 VGND 0.001895f
C1756 VPWR.n104 VGND 0.00196f
C1757 VPWR.n105 VGND 8.22e-19
C1758 VPWR.n106 VGND 8.79e-19
C1759 VPWR.t379 VGND 8.5e-19
C1760 VPWR.t358 VGND 8.5e-19
C1761 VPWR.n107 VGND 0.001889f
C1762 VPWR.n108 VGND 0.004904f
C1763 VPWR.t3 VGND 0.004392f
C1764 VPWR.n109 VGND 0.00508f
C1765 VPWR.t5 VGND 0.001039f
C1766 VPWR.t7 VGND 0.001039f
C1767 VPWR.n110 VGND 0.002121f
C1768 VPWR.n111 VGND 0.001122f
C1769 VPWR.n112 VGND 0.002458f
C1770 VPWR.t459 VGND 8.5e-19
C1771 VPWR.t306 VGND 8.5e-19
C1772 VPWR.n113 VGND 0.001889f
C1773 VPWR.t73 VGND 0.001039f
C1774 VPWR.t1 VGND 0.00141f
C1775 VPWR.n114 VGND 0.002645f
C1776 VPWR.n115 VGND 0.002458f
C1777 VPWR.t132 VGND 0.002797f
C1778 VPWR.t529 VGND 0.005936f
C1779 VPWR.n117 VGND 0.01522f
C1780 VPWR.t133 VGND 0.002797f
C1781 VPWR.n118 VGND 0.00829f
C1782 VPWR.t383 VGND 0.003921f
C1783 VPWR.t489 VGND 0.001447f
C1784 VPWR.t333 VGND 0.001002f
C1785 VPWR.n119 VGND 0.0026f
C1786 VPWR.n120 VGND 0.007599f
C1787 VPWR.n121 VGND 0.004971f
C1788 VPWR.n122 VGND 8.22e-19
C1789 VPWR.t465 VGND 0.00141f
C1790 VPWR.t79 VGND 0.001039f
C1791 VPWR.n123 VGND 0.002645f
C1792 VPWR.n124 VGND 0.001336f
C1793 VPWR.n125 VGND 0.00114f
C1794 VPWR.n126 VGND 0.001639f
C1795 VPWR.n127 VGND 8.79e-19
C1796 VPWR.n128 VGND 0.001099f
C1797 VPWR.n129 VGND 0.00196f
C1798 VPWR.n130 VGND 8.79e-19
C1799 VPWR.n131 VGND 0.001716f
C1800 VPWR.n132 VGND 0.001099f
C1801 VPWR.n133 VGND 8.19e-19
C1802 VPWR.n134 VGND 0.00114f
C1803 VPWR.n135 VGND 0.00483f
C1804 VPWR.n136 VGND 8.2e-19
C1805 VPWR.n137 VGND 4.81e-19
C1806 VPWR.n138 VGND 0.002733f
C1807 VPWR.n139 VGND 0.001122f
C1808 VPWR.n140 VGND 8.2e-19
C1809 VPWR.n141 VGND 0.00483f
C1810 VPWR.n142 VGND 0.004708f
C1811 VPWR.n143 VGND 0.002973f
C1812 VPWR.n144 VGND 7.63e-19
C1813 VPWR.n145 VGND 0.002458f
C1814 VPWR.n146 VGND 0.002084f
C1815 VPWR.n147 VGND 0.001247f
C1816 VPWR.t197 VGND 0.03319f
C1817 VPWR.t341 VGND 0.03382f
C1818 VPWR.t104 VGND 0.009033f
C1819 VPWR.t337 VGND 0.009558f
C1820 VPWR.t339 VGND 0.015755f
C1821 VPWR.t335 VGND 0.007877f
C1822 VPWR.t336 VGND 0.00141f
C1823 VPWR.t375 VGND 0.001039f
C1824 VPWR.n148 VGND 0.002603f
C1825 VPWR.n149 VGND 0.004036f
C1826 VPWR.n150 VGND 0.003278f
C1827 VPWR.t338 VGND 0.001039f
C1828 VPWR.t340 VGND 0.001039f
C1829 VPWR.n151 VGND 0.002108f
C1830 VPWR.t542 VGND 0.011578f
C1831 VPWR.n152 VGND 0.010238f
C1832 VPWR.t198 VGND 0.002797f
C1833 VPWR.t507 VGND 0.005936f
C1834 VPWR.n154 VGND 0.01522f
C1835 VPWR.t199 VGND 0.002797f
C1836 VPWR.n155 VGND 0.00829f
C1837 VPWR.n156 VGND 0.00214f
C1838 VPWR.t206 VGND 0.002797f
C1839 VPWR.t500 VGND 0.005936f
C1840 VPWR.n158 VGND 0.01522f
C1841 VPWR.t207 VGND 0.002797f
C1842 VPWR.n159 VGND 0.00829f
C1843 VPWR.n160 VGND 0.006993f
C1844 VPWR.t342 VGND 0.004348f
C1845 VPWR.n161 VGND 0.005656f
C1846 VPWR.t105 VGND 0.002774f
C1847 VPWR.n162 VGND 0.001098f
C1848 VPWR.n163 VGND 0.003045f
C1849 VPWR.n164 VGND 0.002458f
C1850 VPWR.n165 VGND 0.003278f
C1851 VPWR.n166 VGND 0.006453f
C1852 VPWR.n167 VGND 0.004396f
C1853 VPWR.n168 VGND 0.005733f
C1854 VPWR.t106 VGND 0.002774f
C1855 VPWR.n169 VGND 0.004792f
C1856 VPWR.n170 VGND 0.003242f
C1857 VPWR.n171 VGND 0.001817f
C1858 VPWR.n172 VGND 3.05e-19
C1859 VPWR.n173 VGND 0.001895f
C1860 VPWR.n174 VGND 0.001716f
C1861 VPWR.n175 VGND 0.001099f
C1862 VPWR.n176 VGND 8.19e-19
C1863 VPWR.n177 VGND 7.48e-19
C1864 VPWR.n178 VGND 0.006018f
C1865 VPWR.n179 VGND 0.011793f
C1866 VPWR.t374 VGND 0.011448f
C1867 VPWR.t92 VGND 0.009453f
C1868 VPWR.t86 VGND 0.012814f
C1869 VPWR.t88 VGND 0.018065f
C1870 VPWR.t90 VGND 0.019115f
C1871 VPWR.t359 VGND 0.017015f
C1872 VPWR.t320 VGND 0.022371f
C1873 VPWR.t251 VGND 0.009033f
C1874 VPWR.t314 VGND 0.009558f
C1875 VPWR.t316 VGND 0.018065f
C1876 VPWR.t318 VGND 0.019115f
C1877 VPWR.t58 VGND 0.017015f
C1878 VPWR.t466 VGND 0.019326f
C1879 VPWR.t468 VGND 0.009663f
C1880 VPWR.t462 VGND 0.003256f
C1881 VPWR.t277 VGND 0.009033f
C1882 VPWR.t464 VGND 0.009243f
C1883 VPWR.t427 VGND 0.010083f
C1884 VPWR.t78 VGND 0.01649f
C1885 VPWR.t488 VGND 0.013339f
C1886 VPWR.t332 VGND 0.014284f
C1887 VPWR.t131 VGND 0.008823f
C1888 VPWR.t382 VGND 0.011343f
C1889 VPWR.t72 VGND 0.012919f
C1890 VPWR.t458 VGND 0.010083f
C1891 VPWR.t0 VGND 0.009243f
C1892 VPWR.t305 VGND 0.009033f
C1893 VPWR.t4 VGND 0.006827f
C1894 VPWR.t6 VGND 0.011553f
C1895 VPWR.t2 VGND 0.01691f
C1896 VPWR.t230 VGND 0.036761f
C1897 VPWR.t322 VGND 0.034345f
C1898 VPWR.t328 VGND 0.018065f
C1899 VPWR.t326 VGND 0.018065f
C1900 VPWR.t324 VGND 0.019115f
C1901 VPWR.t287 VGND 0.013444f
C1902 VPWR.t279 VGND 0.01628f
C1903 VPWR.t355 VGND 0.009033f
C1904 VPWR.t285 VGND 0.009243f
C1905 VPWR.t84 VGND 0.009033f
C1906 VPWR.t283 VGND 0.003256f
C1907 VPWR.t281 VGND 0.015965f
C1908 VPWR.t433 VGND 0.011553f
C1909 VPWR.t70 VGND 0.003361f
C1910 VPWR.t66 VGND 0.016175f
C1911 VPWR.t64 VGND 0.010293f
C1912 VPWR.t263 VGND 0.009033f
C1913 VPWR.t68 VGND 0.009033f
C1914 VPWR.t261 VGND 0.010083f
C1915 VPWR.t351 VGND 0.009033f
C1916 VPWR.t259 VGND 0.003361f
C1917 VPWR.t265 VGND 0.015965f
C1918 VPWR.t445 VGND 0.011553f
C1919 VPWR.t347 VGND 0.003361f
C1920 VPWR.t349 VGND 0.016175f
C1921 VPWR.t343 VGND 0.009348f
C1922 VPWR.t399 VGND 0.009033f
C1923 VPWR.t345 VGND 0.009243f
C1924 VPWR.t94 VGND 0.003781f
C1925 VPWR.t401 VGND 0.009663f
C1926 VPWR.t431 VGND 0.01607f
C1927 VPWR.t8 VGND 0.009663f
C1928 VPWR.t357 VGND 0.003256f
C1929 VPWR.t378 VGND 0.009663f
C1930 VPWR.n180 VGND 0.022631f
C1931 VPWR.n181 VGND 0.01224f
C1932 VPWR.n182 VGND 7.7e-19
C1933 VPWR.n183 VGND 0.001122f
C1934 VPWR.n184 VGND 0.001122f
C1935 VPWR.n185 VGND 0.001514f
C1936 VPWR.t9 VGND 8.5e-19
C1937 VPWR.t432 VGND 8.5e-19
C1938 VPWR.n186 VGND 0.001889f
C1939 VPWR.n187 VGND 0.004904f
C1940 VPWR.t402 VGND 0.001039f
C1941 VPWR.t346 VGND 0.00141f
C1942 VPWR.n188 VGND 0.002645f
C1943 VPWR.n189 VGND 0.001122f
C1944 VPWR.n190 VGND 0.001158f
C1945 VPWR.n191 VGND 0.001099f
C1946 VPWR.n192 VGND 0.00196f
C1947 VPWR.n193 VGND 8.79e-19
C1948 VPWR.n194 VGND 0.001099f
C1949 VPWR.n195 VGND 0.001716f
C1950 VPWR.n196 VGND 0.001321f
C1951 VPWR.n197 VGND 0.001817f
C1952 VPWR.t95 VGND 8.5e-19
C1953 VPWR.t400 VGND 8.5e-19
C1954 VPWR.n198 VGND 0.001889f
C1955 VPWR.t344 VGND 0.001039f
C1956 VPWR.t350 VGND 0.001039f
C1957 VPWR.n199 VGND 0.002121f
C1958 VPWR.n200 VGND 0.002458f
C1959 VPWR.t348 VGND 0.004348f
C1960 VPWR.n201 VGND 0.004366f
C1961 VPWR.t446 VGND 0.001039f
C1962 VPWR.t266 VGND 0.00141f
C1963 VPWR.n202 VGND 0.002603f
C1964 VPWR.t260 VGND 0.001039f
C1965 VPWR.t262 VGND 0.001039f
C1966 VPWR.n203 VGND 0.002108f
C1967 VPWR.n204 VGND 0.002292f
C1968 VPWR.n205 VGND 0.003278f
C1969 VPWR.t352 VGND 0.001039f
C1970 VPWR.t69 VGND 0.00141f
C1971 VPWR.n206 VGND 0.002603f
C1972 VPWR.t264 VGND 0.004348f
C1973 VPWR.t65 VGND 0.001039f
C1974 VPWR.t67 VGND 0.001039f
C1975 VPWR.n207 VGND 0.002108f
C1976 VPWR.n208 VGND 0.001098f
C1977 VPWR.t71 VGND 0.004348f
C1978 VPWR.n209 VGND 0.004366f
C1979 VPWR.t434 VGND 0.001039f
C1980 VPWR.t282 VGND 0.00141f
C1981 VPWR.n210 VGND 0.002603f
C1982 VPWR.t85 VGND 8.5e-19
C1983 VPWR.t356 VGND 8.5e-19
C1984 VPWR.n211 VGND 0.001889f
C1985 VPWR.t284 VGND 0.001039f
C1986 VPWR.t286 VGND 0.001039f
C1987 VPWR.n212 VGND 0.002118f
C1988 VPWR.n213 VGND 0.006813f
C1989 VPWR.n214 VGND 9.98e-19
C1990 VPWR.t280 VGND 0.004392f
C1991 VPWR.t288 VGND 0.001039f
C1992 VPWR.t325 VGND 0.00141f
C1993 VPWR.n215 VGND 0.002645f
C1994 VPWR.t361 VGND 0.001039f
C1995 VPWR.t456 VGND 0.00141f
C1996 VPWR.n216 VGND 0.002645f
C1997 VPWR.n217 VGND 0.008525f
C1998 VPWR.n218 VGND 8.19e-19
C1999 VPWR.n219 VGND 0.00114f
C2000 VPWR.n220 VGND 8.79e-19
C2001 VPWR.n221 VGND 0.001099f
C2002 VPWR.n222 VGND 4.3e-19
C2003 VPWR.n223 VGND 0.001099f
C2004 VPWR.n224 VGND 0.0017f
C2005 VPWR.n225 VGND 0.001911f
C2006 VPWR.n226 VGND 0.00196f
C2007 VPWR.n228 VGND 0.001461f
C2008 VPWR.n229 VGND 0.003278f
C2009 VPWR.t327 VGND 0.001039f
C2010 VPWR.t329 VGND 0.001039f
C2011 VPWR.n230 VGND 0.002121f
C2012 VPWR.t453 VGND 0.001039f
C2013 VPWR.t454 VGND 0.001039f
C2014 VPWR.n231 VGND 0.002121f
C2015 VPWR.t323 VGND 0.004392f
C2016 VPWR.t455 VGND 0.004392f
C2017 VPWR.n232 VGND 0.008822f
C2018 VPWR.t231 VGND 0.002797f
C2019 VPWR.t495 VGND 0.005936f
C2020 VPWR.n234 VGND 0.01522f
C2021 VPWR.t232 VGND 0.002797f
C2022 VPWR.n235 VGND 0.00829f
C2023 VPWR.t247 VGND 0.002797f
C2024 VPWR.t538 VGND 0.005936f
C2025 VPWR.n237 VGND 0.01522f
C2026 VPWR.t248 VGND 0.002797f
C2027 VPWR.n238 VGND 0.00829f
C2028 VPWR.n239 VGND 0.006895f
C2029 VPWR.n240 VGND 0.002757f
C2030 VPWR.n241 VGND 0.002458f
C2031 VPWR.n242 VGND 0.003278f
C2032 VPWR.n243 VGND 7.63e-19
C2033 VPWR.n244 VGND 0.004881f
C2034 VPWR.n245 VGND 7.57e-19
C2035 VPWR.n246 VGND 0.001817f
C2036 VPWR.n247 VGND 0.001321f
C2037 VPWR.n248 VGND 0.0017f
C2038 VPWR.n249 VGND 0.001911f
C2039 VPWR.n250 VGND 0.00196f
C2040 VPWR.n251 VGND 8.79e-19
C2041 VPWR.n252 VGND 0.001099f
C2042 VPWR.n253 VGND 0.001336f
C2043 VPWR.n254 VGND 6.24e-19
C2044 VPWR.n255 VGND 8.9e-19
C2045 VPWR.n256 VGND 0.005263f
C2046 VPWR.n257 VGND 7.07e-19
C2047 VPWR.n258 VGND 0.002458f
C2048 VPWR.n259 VGND 0.002975f
C2049 VPWR.n260 VGND 0.001122f
C2050 VPWR.n261 VGND 9.15e-19
C2051 VPWR.n262 VGND 0.004109f
C2052 VPWR.n263 VGND 1.01e-19
C2053 VPWR.n264 VGND 0.002156f
C2054 VPWR.n265 VGND 0.001122f
C2055 VPWR.n266 VGND 0.002458f
C2056 VPWR.n267 VGND 5.87e-19
C2057 VPWR.n268 VGND 0.001775f
C2058 VPWR.n269 VGND 0.00436f
C2059 VPWR.n270 VGND 0.00106f
C2060 VPWR.n271 VGND 0.004109f
C2061 VPWR.n272 VGND 4.42e-20
C2062 VPWR.n273 VGND 0.002975f
C2063 VPWR.n274 VGND 0.001122f
C2064 VPWR.n275 VGND 0.001117f
C2065 VPWR.n276 VGND 0.004109f
C2066 VPWR.n277 VGND 1.01e-19
C2067 VPWR.n278 VGND 0.002156f
C2068 VPWR.n279 VGND 0.001122f
C2069 VPWR.n280 VGND 9.46e-19
C2070 VPWR.n281 VGND 0.002973f
C2071 VPWR.n282 VGND 0.004708f
C2072 VPWR.n283 VGND 0.00483f
C2073 VPWR.n284 VGND 7.95e-19
C2074 VPWR.n285 VGND 6.24e-19
C2075 VPWR.n286 VGND 8.19e-19
C2076 VPWR.n287 VGND 0.001099f
C2077 VPWR.n288 VGND 0.001716f
C2078 VPWR.n289 VGND 0.001895f
C2079 VPWR.n290 VGND 0.105698f
C2080 VPWR.n291 VGND 0.001895f
C2081 VPWR.n292 VGND 0.00196f
C2082 VPWR.n293 VGND 3.05e-19
C2083 VPWR.n294 VGND 0.001716f
C2084 VPWR.n295 VGND 5.17e-19
C2085 VPWR.n296 VGND 0.001099f
C2086 VPWR.n297 VGND 0.00196f
C2087 VPWR.n298 VGND 8.79e-19
C2088 VPWR.n299 VGND 0.001318f
C2089 VPWR.n300 VGND 0.001099f
C2090 VPWR.n301 VGND 8.79e-19
C2091 VPWR.n302 VGND 8.19e-19
C2092 VPWR.n303 VGND 0.001099f
C2093 VPWR.n304 VGND 0.001716f
C2094 VPWR.n305 VGND 0.001895f
C2095 VPWR.n306 VGND 0.129213f
C2096 VPWR.n307 VGND 0.129213f
C2097 VPWR.n308 VGND 0.00196f
C2098 VPWR.n309 VGND 0.002458f
C2099 VPWR.t543 VGND 0.016311f
C2100 VPWR.t522 VGND 0.040428f
C2101 VPWR.n310 VGND 0.018883f
C2102 VPWR.t122 VGND 0.028988f
C2103 VPWR.t407 VGND 0.011448f
C2104 VPWR.t145 VGND 0.009033f
C2105 VPWR.t405 VGND 0.014389f
C2106 VPWR.t403 VGND 0.012184f
C2107 VPWR.t409 VGND 0.012288f
C2108 VPWR.t10 VGND 0.010083f
C2109 VPWR.t82 VGND 0.007037f
C2110 VPWR.t393 VGND 0.009663f
C2111 VPWR.t307 VGND 0.011133f
C2112 VPWR.t478 VGND 0.028043f
C2113 VPWR.t472 VGND 0.015649f
C2114 VPWR.t447 VGND 0.01859f
C2115 VPWR.t396 VGND 0.010293f
C2116 VPWR.t222 VGND 0.009978f
C2117 VPWR.t11 VGND 0.022371f
C2118 VPWR.t62 VGND 0.01607f
C2119 VPWR.t56 VGND 0.022161f
C2120 VPWR.t225 VGND 0.045268f
C2121 VPWR.t157 VGND 0.032244f
C2122 VPWR.n311 VGND 0.020826f
C2123 VPWR.t215 VGND 0.003052f
C2124 VPWR.n312 VGND 0.003857f
C2125 VPWR.n313 VGND 0.002975f
C2126 VPWR.t162 VGND 0.003052f
C2127 VPWR.n314 VGND 0.003857f
C2128 VPWR.n315 VGND 0.003278f
C2129 VPWR.n316 VGND 0.005211f
C2130 VPWR.n317 VGND 0.001817f
C2131 VPWR.t521 VGND 0.040428f
C2132 VPWR.n318 VGND 0.020138f
C2133 VPWR.n319 VGND 0.001639f
C2134 VPWR.n320 VGND 0.001321f
C2135 VPWR.n321 VGND 8.79e-19
C2136 VPWR.n322 VGND 0.001099f
C2137 VPWR.n323 VGND 8.79e-19
C2138 VPWR.n324 VGND 3.05e-19
C2139 VPWR.t112 VGND 0.003052f
C2140 VPWR.n325 VGND 0.003857f
C2141 VPWR.n326 VGND 0.002975f
C2142 VPWR.t184 VGND 0.003052f
C2143 VPWR.n327 VGND 0.003857f
C2144 VPWR.n328 VGND 0.003278f
C2145 VPWR.n329 VGND 0.005211f
C2146 VPWR.n330 VGND 0.003278f
C2147 VPWR.t515 VGND 0.040428f
C2148 VPWR.n331 VGND 0.020138f
C2149 VPWR.t183 VGND 0.003062f
C2150 VPWR.n332 VGND 8.47e-19
C2151 VPWR.t165 VGND 0.002815f
C2152 VPWR.n333 VGND 0.004233f
C2153 VPWR.n334 VGND 0.002814f
C2154 VPWR.n335 VGND 8.79e-19
C2155 VPWR.n336 VGND 0.00196f
C2156 VPWR.n337 VGND 0.001895f
C2157 VPWR.n338 VGND 0.00196f
C2158 VPWR.n339 VGND 0.001798f
C2159 VPWR.n340 VGND 8.79e-19
C2160 VPWR.t188 VGND 0.038756f
C2161 VPWR.t98 VGND 0.019221f
C2162 VPWR.t330 VGND 0.007877f
C2163 VPWR.t474 VGND 0.009663f
C2164 VPWR.t391 VGND 0.01628f
C2165 VPWR.t179 VGND 0.008823f
C2166 VPWR.t440 VGND 0.013864f
C2167 VPWR.t52 VGND 0.019956f
C2168 VPWR.t54 VGND 0.019746f
C2169 VPWR.t484 VGND 0.01901f
C2170 VPWR.t387 VGND 0.020061f
C2171 VPWR.t38 VGND 0.026363f
C2172 VPWR.t191 VGND 0.01817f
C2173 VPWR.t385 VGND 0.019746f
C2174 VPWR.t470 VGND 0.01901f
C2175 VPWR.t299 VGND 0.020061f
C2176 VPWR.t380 VGND 0.029409f
C2177 VPWR.t185 VGND 0.054931f
C2178 VPWR.t244 VGND 0.041907f
C2179 VPWR.n341 VGND 0.020826f
C2180 VPWR.t100 VGND 0.002816f
C2181 VPWR.n342 VGND 0.002713f
C2182 VPWR.n343 VGND 0.011617f
C2183 VPWR.t545 VGND 0.011732f
C2184 VPWR.n344 VGND 0.012856f
C2185 VPWR.t99 VGND 0.002774f
C2186 VPWR.n345 VGND 0.004047f
C2187 VPWR.n346 VGND 0.003991f
C2188 VPWR.t189 VGND 0.002797f
C2189 VPWR.t509 VGND 0.005936f
C2190 VPWR.n348 VGND 0.01522f
C2191 VPWR.t190 VGND 0.002797f
C2192 VPWR.n349 VGND 0.00829f
C2193 VPWR.t249 VGND 0.002797f
C2194 VPWR.t537 VGND 0.005936f
C2195 VPWR.n351 VGND 0.01522f
C2196 VPWR.t250 VGND 0.002797f
C2197 VPWR.n352 VGND 0.00829f
C2198 VPWR.n353 VGND 0.00683f
C2199 VPWR.n354 VGND 0.00214f
C2200 VPWR.n355 VGND 0.001961f
C2201 VPWR.n356 VGND 0.001552f
C2202 VPWR.n357 VGND 0.003924f
C2203 VPWR.t245 VGND 0.003062f
C2204 VPWR.n358 VGND 0.006245f
C2205 VPWR.t539 VGND 0.040639f
C2206 VPWR.n359 VGND 0.018085f
C2207 VPWR.n360 VGND 0.001099f
C2208 VPWR.n361 VGND 0.00196f
C2209 VPWR.n362 VGND 8.79e-19
C2210 VPWR.n363 VGND 0.003278f
C2211 VPWR.t510 VGND 0.020527f
C2212 VPWR.n364 VGND 0.011575f
C2213 VPWR.n365 VGND 0.003278f
C2214 VPWR.t246 VGND 0.003052f
C2215 VPWR.t187 VGND 0.002774f
C2216 VPWR.n366 VGND 0.006677f
C2217 VPWR.t192 VGND 0.003052f
C2218 VPWR.n367 VGND 0.002371f
C2219 VPWR.n368 VGND 0.003278f
C2220 VPWR.t381 VGND 0.00141f
C2221 VPWR.t300 VGND 0.001447f
C2222 VPWR.n369 VGND 0.00301f
C2223 VPWR.t502 VGND 0.040428f
C2224 VPWR.n370 VGND 0.018233f
C2225 VPWR.n371 VGND 0.001817f
C2226 VPWR.t386 VGND 6.35e-19
C2227 VPWR.t471 VGND 0.001025f
C2228 VPWR.n372 VGND 0.003075f
C2229 VPWR.n373 VGND 0.004788f
C2230 VPWR.n374 VGND 0.002717f
C2231 VPWR.n375 VGND 0.003278f
C2232 VPWR.n376 VGND 0.003278f
C2233 VPWR.n377 VGND 0.003166f
C2234 VPWR.n378 VGND 0.002784f
C2235 VPWR.n379 VGND 0.005297f
C2236 VPWR.n380 VGND 0.003278f
C2237 VPWR.n381 VGND 0.003278f
C2238 VPWR.n382 VGND 0.002458f
C2239 VPWR.n383 VGND 0.001597f
C2240 VPWR.n384 VGND 0.004263f
C2241 VPWR.n385 VGND 0.001942f
C2242 VPWR.n386 VGND 0.003278f
C2243 VPWR.n387 VGND 0.011197f
C2244 VPWR.n388 VGND 0.011575f
C2245 VPWR.n389 VGND 0.011575f
C2246 VPWR.n390 VGND 0.003278f
C2247 VPWR.n391 VGND 0.003278f
C2248 VPWR.n392 VGND 0.003278f
C2249 VPWR.n393 VGND 0.008555f
C2250 VPWR.n394 VGND 0.029171f
C2251 VPWR.n395 VGND 0.00843f
C2252 VPWR.t186 VGND 0.002774f
C2253 VPWR.n396 VGND 0.006371f
C2254 VPWR.n397 VGND 0.004028f
C2255 VPWR.n398 VGND 0.001817f
C2256 VPWR.n399 VGND 8.22e-19
C2257 VPWR.n400 VGND 0.001716f
C2258 VPWR.n401 VGND 0.001099f
C2259 VPWR.n402 VGND 4.28e-19
C2260 VPWR.n403 VGND 0.00114f
C2261 VPWR.n404 VGND 0.003413f
C2262 VPWR.n405 VGND 0.008994f
C2263 VPWR.n406 VGND 7.48e-19
C2264 VPWR.n407 VGND 8.19e-19
C2265 VPWR.n408 VGND 0.001099f
C2266 VPWR.n409 VGND 0.001716f
C2267 VPWR.n410 VGND 0.001895f
C2268 VPWR.n411 VGND 0.129213f
C2269 VPWR.n412 VGND 0.001895f
C2270 VPWR.n413 VGND 0.09976f
C2271 VPWR.n414 VGND 0.00196f
C2272 VPWR.n415 VGND 0.004028f
C2273 VPWR.n416 VGND 8.79e-19
C2274 VPWR.t126 VGND 0.002797f
C2275 VPWR.t534 VGND 0.005936f
C2276 VPWR.n418 VGND 0.01522f
C2277 VPWR.t127 VGND 0.002797f
C2278 VPWR.n419 VGND 0.00829f
C2279 VPWR.t177 VGND 0.002797f
C2280 VPWR.t505 VGND 0.005936f
C2281 VPWR.n421 VGND 0.01522f
C2282 VPWR.t178 VGND 0.002797f
C2283 VPWR.n422 VGND 0.00829f
C2284 VPWR.n423 VGND 0.00683f
C2285 VPWR.t508 VGND 0.011578f
C2286 VPWR.t201 VGND 0.002804f
C2287 VPWR.n424 VGND 0.016794f
C2288 VPWR.t202 VGND 0.002945f
C2289 VPWR.n425 VGND 0.018712f
C2290 VPWR.n426 VGND 0.00214f
C2291 VPWR.n427 VGND 0.003649f
C2292 VPWR.n428 VGND 0.006048f
C2293 VPWR.n429 VGND 0.007142f
C2294 VPWR.t499 VGND 0.020814f
C2295 VPWR.t211 VGND 0.002774f
C2296 VPWR.n430 VGND 0.034853f
C2297 VPWR.n431 VGND 0.009157f
C2298 VPWR.n432 VGND 0.008604f
C2299 VPWR.t125 VGND 0.041697f
C2300 VPWR.t200 VGND 0.050099f
C2301 VPWR.t210 VGND 0.007877f
C2302 VPWR.t311 VGND 0.003512f
C2303 VPWR.n433 VGND 0.004071f
C2304 VPWR.n434 VGND 0.003278f
C2305 VPWR.n435 VGND 0.007102f
C2306 VPWR.n436 VGND 0.003278f
C2307 VPWR.t536 VGND 0.040428f
C2308 VPWR.n437 VGND 0.020369f
C2309 VPWR.n438 VGND 0.001817f
C2310 VPWR.t541 VGND 0.040428f
C2311 VPWR.t255 VGND 0.003052f
C2312 VPWR.n439 VGND 0.003857f
C2313 VPWR.n440 VGND 0.001639f
C2314 VPWR.n441 VGND 0.001321f
C2315 VPWR.n442 VGND 8.79e-19
C2316 VPWR.n443 VGND 0.00196f
C2317 VPWR.n445 VGND 0.001911f
C2318 VPWR.n446 VGND 0.00196f
C2319 VPWR.n447 VGND 0.001099f
C2320 VPWR.n448 VGND 0.001461f
C2321 VPWR.n449 VGND 0.001942f
C2322 VPWR.n450 VGND 0.007102f
C2323 VPWR.t208 VGND 0.003064f
C2324 VPWR.n451 VGND 0.003453f
C2325 VPWR.t304 VGND 8.5e-19
C2326 VPWR.t61 VGND 8.5e-19
C2327 VPWR.n452 VGND 0.001849f
C2328 VPWR.n453 VGND 0.003166f
C2329 VPWR.n454 VGND 0.003278f
C2330 VPWR.t497 VGND 0.040428f
C2331 VPWR.n455 VGND 0.018883f
C2332 VPWR.t518 VGND 0.011578f
C2333 VPWR.t143 VGND 0.002804f
C2334 VPWR.n456 VGND 0.016794f
C2335 VPWR.t144 VGND 0.002945f
C2336 VPWR.n457 VGND 0.004131f
C2337 VPWR.t169 VGND 0.028988f
C2338 VPWR.t40 VGND 0.012499f
C2339 VPWR.t411 VGND 0.009453f
C2340 VPWR.t241 VGND 0.01628f
C2341 VPWR.n458 VGND 0.002092f
C2342 VPWR.n459 VGND 7.48e-19
C2343 VPWR.t243 VGND 0.002774f
C2344 VPWR.n460 VGND 0.004886f
C2345 VPWR.n461 VGND 0.002975f
C2346 VPWR.t41 VGND 8.5e-19
C2347 VPWR.t412 VGND 8.5e-19
C2348 VPWR.n462 VGND 0.001849f
C2349 VPWR.t540 VGND 0.011578f
C2350 VPWR.t170 VGND 0.002797f
C2351 VPWR.t504 VGND 0.005936f
C2352 VPWR.n464 VGND 0.01522f
C2353 VPWR.t171 VGND 0.002797f
C2354 VPWR.n465 VGND 0.00829f
C2355 VPWR.t220 VGND 0.002797f
C2356 VPWR.t492 VGND 0.005936f
C2357 VPWR.n467 VGND 0.01522f
C2358 VPWR.t221 VGND 0.002797f
C2359 VPWR.n468 VGND 0.00829f
C2360 VPWR.n469 VGND 0.006993f
C2361 VPWR.n470 VGND 0.00214f
C2362 VPWR.n471 VGND 0.001122f
C2363 VPWR.n472 VGND 0.003045f
C2364 VPWR.t242 VGND 0.002774f
C2365 VPWR.n473 VGND 0.002735f
C2366 VPWR.n474 VGND 0.010472f
C2367 VPWR.n475 VGND 0.010028f
C2368 VPWR.n476 VGND 0.008324f
C2369 VPWR.n477 VGND 0.002458f
C2370 VPWR.n478 VGND 8.19e-19
C2371 VPWR.n479 VGND 0.001099f
C2372 VPWR.n480 VGND 8.79e-19
C2373 VPWR.n481 VGND 8.79e-19
C2374 VPWR.n482 VGND 0.001099f
C2375 VPWR.n483 VGND 0.001099f
C2376 VPWR.n484 VGND 0.00114f
C2377 VPWR.n485 VGND 4.28e-19
C2378 VPWR.n486 VGND 0.003278f
C2379 VPWR.n487 VGND 0.004271f
C2380 VPWR.t524 VGND 0.016311f
C2381 VPWR.n488 VGND 0.002166f
C2382 VPWR.t137 VGND 0.002774f
C2383 VPWR.n489 VGND 0.005961f
C2384 VPWR.t523 VGND 0.019764f
C2385 VPWR.n490 VGND 0.013953f
C2386 VPWR.n491 VGND 0.016048f
C2387 VPWR.n492 VGND 0.001942f
C2388 VPWR.t102 VGND 0.003064f
C2389 VPWR.n493 VGND 0.003417f
C2390 VPWR.n494 VGND 0.003278f
C2391 VPWR.t530 VGND 0.040428f
C2392 VPWR.n495 VGND 0.020369f
C2393 VPWR.n496 VGND 0.003278f
C2394 VPWR.t547 VGND 0.040428f
C2395 VPWR.n497 VGND 0.007102f
C2396 VPWR.n498 VGND 0.001461f
C2397 VPWR.n499 VGND 8.79e-19
C2398 VPWR.n500 VGND 0.007102f
C2399 VPWR.n501 VGND 0.00114f
C2400 VPWR.n502 VGND 0.00114f
C2401 VPWR.n503 VGND 0.001639f
C2402 VPWR.n504 VGND 0.001099f
C2403 VPWR.n505 VGND 0.00196f
C2404 VPWR.n506 VGND 8.79e-19
C2405 VPWR.n507 VGND 0.001099f
C2406 VPWR.n508 VGND 0.0017f
C2407 VPWR.n509 VGND 0.001321f
C2408 VPWR.n510 VGND 0.001817f
C2409 VPWR.n511 VGND 0.003278f
C2410 VPWR.n512 VGND 0.007102f
C2411 VPWR.n513 VGND 0.005211f
C2412 VPWR.n514 VGND 0.020369f
C2413 VPWR.n515 VGND 0.003551f
C2414 VPWR.n516 VGND 0.003278f
C2415 VPWR.n517 VGND 0.003278f
C2416 VPWR.n518 VGND 0.005442f
C2417 VPWR.n519 VGND 0.00687f
C2418 VPWR.t234 VGND 0.003052f
C2419 VPWR.n520 VGND 0.003857f
C2420 VPWR.n521 VGND 0.002586f
C2421 VPWR.n522 VGND 0.002458f
C2422 VPWR.n523 VGND 0.001122f
C2423 VPWR.n524 VGND 0.001523f
C2424 VPWR.t138 VGND 0.002819f
C2425 VPWR.n525 VGND 0.003761f
C2426 VPWR.n526 VGND 0.009536f
C2427 VPWR.t115 VGND 0.002774f
C2428 VPWR.n527 VGND 0.008608f
C2429 VPWR.n528 VGND 0.015524f
C2430 VPWR.n529 VGND 0.003278f
C2431 VPWR.n530 VGND 0.003278f
C2432 VPWR.n531 VGND 0.003278f
C2433 VPWR.n532 VGND 0.015873f
C2434 VPWR.n533 VGND 0.015659f
C2435 VPWR.n534 VGND 0.021492f
C2436 VPWR.t114 VGND 0.002774f
C2437 VPWR.n535 VGND 0.008608f
C2438 VPWR.n536 VGND 0.003053f
C2439 VPWR.n537 VGND 0.001817f
C2440 VPWR.n538 VGND 8.22e-19
C2441 VPWR.n539 VGND 0.001716f
C2442 VPWR.n540 VGND 0.001895f
C2443 VPWR.n541 VGND 0.00196f
C2444 VPWR.n542 VGND 0.00196f
C2445 VPWR.n543 VGND 0.001895f
C2446 VPWR.n544 VGND 0.001716f
C2447 VPWR.n545 VGND 3.05e-19
C2448 VPWR.n546 VGND 9.98e-19
C2449 VPWR.n547 VGND 0.003045f
C2450 VPWR.n548 VGND 0.01215f
C2451 VPWR.n549 VGND 0.022736f
C2452 VPWR.t113 VGND 0.058187f
C2453 VPWR.t101 VGND 0.061023f
C2454 VPWR.t233 VGND 0.054931f
C2455 VPWR.t303 VGND 0.012499f
C2456 VPWR.t60 VGND 0.038441f
C2457 VPWR.t142 VGND 0.045478f
C2458 VPWR.t107 VGND 0.036761f
C2459 VPWR.t295 VGND 0.034345f
C2460 VPWR.t293 VGND 0.018065f
C2461 VPWR.t291 VGND 0.018065f
C2462 VPWR.t297 VGND 0.019115f
C2463 VPWR.t376 VGND 0.013444f
C2464 VPWR.t384 VGND 0.006827f
C2465 VPWR.t76 VGND 0.008823f
C2466 VPWR.t442 VGND 0.010083f
C2467 VPWR.t273 VGND 0.008823f
C2468 VPWR.t486 VGND 0.009033f
C2469 VPWR.t271 VGND 0.010608f
C2470 VPWR.t269 VGND 0.012604f
C2471 VPWR.t275 VGND 0.019326f
C2472 VPWR.t74 VGND 0.01607f
C2473 VPWR.t257 VGND 0.022161f
C2474 VPWR.t148 VGND 0.035605f
C2475 VPWR.t203 VGND 0.061023f
C2476 VPWR.n550 VGND 0.030803f
C2477 VPWR.n551 VGND 0.00348f
C2478 VPWR.n552 VGND 3.05e-19
C2479 VPWR.t209 VGND 0.003064f
C2480 VPWR.n553 VGND 0.003485f
C2481 VPWR.n554 VGND 0.005678f
C2482 VPWR.t501 VGND 0.019759f
C2483 VPWR.t149 VGND 0.003052f
C2484 VPWR.n555 VGND 0.006093f
C2485 VPWR.n556 VGND 0.005599f
C2486 VPWR.n557 VGND 0.00887f
C2487 VPWR.n558 VGND 0.001461f
C2488 VPWR.n559 VGND 0.001099f
C2489 VPWR.n560 VGND 0.00196f
C2490 VPWR.n561 VGND 0.00196f
C2491 VPWR.n562 VGND 8.79e-19
C2492 VPWR.n563 VGND 0.00114f
C2493 VPWR.n564 VGND 8.79e-19
C2494 VPWR.n565 VGND 0.001099f
C2495 VPWR.n566 VGND 0.001639f
C2496 VPWR.n567 VGND 0.00114f
C2497 VPWR.n568 VGND 0.001336f
C2498 VPWR.n569 VGND 0.001099f
C2499 VPWR.n570 VGND 0.001716f
C2500 VPWR.n571 VGND 0.001895f
C2501 VPWR.n572 VGND 0.09976f
C2502 VPWR.n573 VGND 0.001895f
C2503 VPWR.n574 VGND 0.001716f
C2504 VPWR.n575 VGND 0.001321f
C2505 VPWR.n576 VGND 0.003278f
C2506 VPWR.t513 VGND 0.040428f
C2507 VPWR.n577 VGND 0.022605f
C2508 VPWR.n578 VGND 0.003937f
C2509 VPWR.n579 VGND 0.002458f
C2510 VPWR.t258 VGND 8.5e-19
C2511 VPWR.t75 VGND 8.5e-19
C2512 VPWR.n580 VGND 0.001849f
C2513 VPWR.t276 VGND 0.004348f
C2514 VPWR.n581 VGND 0.005716f
C2515 VPWR.t150 VGND 0.003052f
C2516 VPWR.n582 VGND 0.002124f
C2517 VPWR.t487 VGND 0.003815f
C2518 VPWR.n583 VGND 0.002975f
C2519 VPWR.t270 VGND 0.001039f
C2520 VPWR.t272 VGND 0.001039f
C2521 VPWR.n584 VGND 0.002118f
C2522 VPWR.t274 VGND 0.00141f
C2523 VPWR.t77 VGND 0.001039f
C2524 VPWR.n585 VGND 0.002645f
C2525 VPWR.n586 VGND 0.005038f
C2526 VPWR.n587 VGND 2.87e-19
C2527 VPWR.t377 VGND 0.001039f
C2528 VPWR.t438 VGND 0.00141f
C2529 VPWR.n588 VGND 0.002645f
C2530 VPWR.t457 VGND 0.001039f
C2531 VPWR.t298 VGND 0.00141f
C2532 VPWR.n589 VGND 0.002645f
C2533 VPWR.n590 VGND 0.008525f
C2534 VPWR.n591 VGND 8.19e-19
C2535 VPWR.n592 VGND 0.00114f
C2536 VPWR.n593 VGND 8.79e-19
C2537 VPWR.n594 VGND 0.001099f
C2538 VPWR.n595 VGND 0.00196f
C2539 VPWR.n596 VGND 0.001099f
C2540 VPWR.n597 VGND 0.001716f
C2541 VPWR.n598 VGND 0.001895f
C2542 VPWR.n599 VGND 0.09976f
C2543 VPWR.n600 VGND 0.001461f
C2544 VPWR.n601 VGND 0.003278f
C2545 VPWR.t435 VGND 0.001039f
C2546 VPWR.t436 VGND 0.001039f
C2547 VPWR.n602 VGND 0.002121f
C2548 VPWR.t292 VGND 0.001039f
C2549 VPWR.t294 VGND 0.001039f
C2550 VPWR.n603 VGND 0.002121f
C2551 VPWR.t437 VGND 0.004392f
C2552 VPWR.t296 VGND 0.004392f
C2553 VPWR.n604 VGND 0.008822f
C2554 VPWR.t216 VGND 0.002797f
C2555 VPWR.t491 VGND 0.005936f
C2556 VPWR.n606 VGND 0.01522f
C2557 VPWR.t217 VGND 0.002797f
C2558 VPWR.n607 VGND 0.00829f
C2559 VPWR.t108 VGND 0.002797f
C2560 VPWR.t532 VGND 0.005936f
C2561 VPWR.n609 VGND 0.01522f
C2562 VPWR.t109 VGND 0.002797f
C2563 VPWR.n610 VGND 0.00829f
C2564 VPWR.n611 VGND 0.006895f
C2565 VPWR.n612 VGND 0.002757f
C2566 VPWR.n613 VGND 0.002458f
C2567 VPWR.n614 VGND 0.003278f
C2568 VPWR.n615 VGND 7.63e-19
C2569 VPWR.n616 VGND 0.004881f
C2570 VPWR.n617 VGND 7.57e-19
C2571 VPWR.n618 VGND 0.001817f
C2572 VPWR.n619 VGND 0.001321f
C2573 VPWR.n620 VGND 0.001716f
C2574 VPWR.n621 VGND 0.001895f
C2575 VPWR.n622 VGND 0.00196f
C2576 VPWR.n623 VGND 8.79e-19
C2577 VPWR.n624 VGND 0.001099f
C2578 VPWR.n625 VGND 0.001336f
C2579 VPWR.n626 VGND 6.24e-19
C2580 VPWR.n627 VGND 0.001003f
C2581 VPWR.n628 VGND 0.001003f
C2582 VPWR.n629 VGND 0.001817f
C2583 VPWR.n630 VGND 0.003278f
C2584 VPWR.n631 VGND 0.003278f
C2585 VPWR.n632 VGND 7.07e-19
C2586 VPWR.n633 VGND 0.007026f
C2587 VPWR.n634 VGND 0.001493f
C2588 VPWR.n635 VGND 0.001942f
C2589 VPWR.n636 VGND 0.002458f
C2590 VPWR.n637 VGND 0.001931f
C2591 VPWR.n638 VGND 0.002447f
C2592 VPWR.n639 VGND 0.007706f
C2593 VPWR.n640 VGND 0.003278f
C2594 VPWR.n641 VGND 0.002458f
C2595 VPWR.n642 VGND 0.001942f
C2596 VPWR.n643 VGND 0.004983f
C2597 VPWR.t205 VGND 0.002774f
C2598 VPWR.n644 VGND 0.006371f
C2599 VPWR.n645 VGND 0.011197f
C2600 VPWR.n646 VGND 0.008492f
C2601 VPWR.n647 VGND 0.003278f
C2602 VPWR.n648 VGND 0.003278f
C2603 VPWR.n649 VGND 0.001817f
C2604 VPWR.n650 VGND 0.011386f
C2605 VPWR.n651 VGND 0.013393f
C2606 VPWR.n652 VGND 0.013647f
C2607 VPWR.n653 VGND 0.007161f
C2608 VPWR.t204 VGND 0.002794f
C2609 VPWR.n654 VGND 0.001298f
C2610 VPWR.n655 VGND 0.002021f
C2611 VPWR.n656 VGND 9.98e-19
C2612 VPWR.n657 VGND 0.002084f
C2613 VPWR.n658 VGND 0.002458f
C2614 VPWR.n659 VGND 0.004131f
C2615 VPWR.n660 VGND 0.009645f
C2616 VPWR.n661 VGND 0.001247f
C2617 VPWR.n662 VGND 0.001942f
C2618 VPWR.n663 VGND 0.003278f
C2619 VPWR.n664 VGND 0.003099f
C2620 VPWR.n665 VGND 0.019712f
C2621 VPWR.n666 VGND 0.003099f
C2622 VPWR.n667 VGND 0.003031f
C2623 VPWR.n668 VGND 0.002458f
C2624 VPWR.n669 VGND 0.002458f
C2625 VPWR.n670 VGND 0.002975f
C2626 VPWR.n671 VGND 0.007706f
C2627 VPWR.n672 VGND 0.00348f
C2628 VPWR.n673 VGND 0.001639f
C2629 VPWR.n674 VGND 0.001639f
C2630 VPWR.n675 VGND 9.2e-19
C2631 VPWR.t235 VGND 0.003063f
C2632 VPWR.n676 VGND 0.003435f
C2633 VPWR.n677 VGND 0.002636f
C2634 VPWR.t103 VGND 0.003052f
C2635 VPWR.n678 VGND 0.003857f
C2636 VPWR.n679 VGND 0.00687f
C2637 VPWR.n680 VGND 0.001817f
C2638 VPWR.n681 VGND 0.001321f
C2639 VPWR.n682 VGND 0.0017f
C2640 VPWR.n683 VGND 0.001911f
C2641 VPWR.n684 VGND 0.09976f
C2642 VPWR.n685 VGND 0.00196f
C2643 VPWR.n686 VGND 3.05e-19
C2644 VPWR.n687 VGND 0.001099f
C2645 VPWR.n688 VGND 8.79e-19
C2646 VPWR.t120 VGND 0.003064f
C2647 VPWR.t156 VGND 0.003063f
C2648 VPWR.n689 VGND 0.003435f
C2649 VPWR.n690 VGND 0.003278f
C2650 VPWR.n691 VGND 0.007102f
C2651 VPWR.n692 VGND 0.003278f
C2652 VPWR.t514 VGND 0.040428f
C2653 VPWR.n693 VGND 0.020369f
C2654 VPWR.n694 VGND 0.003278f
C2655 VPWR.t516 VGND 0.040428f
C2656 VPWR.t155 VGND 0.003052f
C2657 VPWR.n695 VGND 0.003857f
C2658 VPWR.t175 VGND 0.003064f
C2659 VPWR.t212 VGND 0.002819f
C2660 VPWR.n696 VGND 0.004155f
C2661 VPWR.n697 VGND 0.001461f
C2662 VPWR.n698 VGND 0.00114f
C2663 VPWR.n699 VGND 0.001099f
C2664 VPWR.n700 VGND 0.00196f
C2665 VPWR.n701 VGND 8.79e-19
C2666 VPWR.n702 VGND 0.001099f
C2667 VPWR.n703 VGND 0.001716f
C2668 VPWR.n704 VGND 0.001321f
C2669 VPWR.n705 VGND 0.010574f
C2670 VPWR.n706 VGND 6.24e-19
C2671 VPWR.n707 VGND 0.001122f
C2672 VPWR.n708 VGND 0.001523f
C2673 VPWR.n709 VGND 0.003417f
C2674 VPWR.n710 VGND 0.002586f
C2675 VPWR.n711 VGND 0.002458f
C2676 VPWR.n712 VGND 0.003278f
C2677 VPWR.n713 VGND 0.00687f
C2678 VPWR.n714 VGND 0.005442f
C2679 VPWR.n715 VGND 0.020369f
C2680 VPWR.n716 VGND 0.003551f
C2681 VPWR.n717 VGND 0.003278f
C2682 VPWR.n718 VGND 0.003278f
C2683 VPWR.n719 VGND 0.005211f
C2684 VPWR.n720 VGND 0.007102f
C2685 VPWR.n721 VGND 0.007102f
C2686 VPWR.n722 VGND 0.003278f
C2687 VPWR.n723 VGND 0.003278f
C2688 VPWR.n724 VGND 0.003278f
C2689 VPWR.n725 VGND 0.007102f
C2690 VPWR.n726 VGND 0.00687f
C2691 VPWR.t176 VGND 0.003052f
C2692 VPWR.n727 VGND 0.003857f
C2693 VPWR.n728 VGND 0.002636f
C2694 VPWR.n729 VGND 0.001942f
C2695 VPWR.n730 VGND 0.001514f
C2696 VPWR.n731 VGND 9.2e-19
C2697 VPWR.n732 VGND 0.003417f
C2698 VPWR.n733 VGND 0.002586f
C2699 VPWR.n734 VGND 0.00114f
C2700 VPWR.n735 VGND 0.001336f
C2701 VPWR.n736 VGND 0.001099f
C2702 VPWR.n737 VGND 0.001716f
C2703 VPWR.n738 VGND 0.001895f
C2704 VPWR.n739 VGND 0.129213f
C2705 VPWR.n740 VGND 0.001895f
C2706 VPWR.n741 VGND 0.001716f
C2707 VPWR.n742 VGND 0.001099f
C2708 VPWR.n743 VGND 0.001461f
C2709 VPWR.n744 VGND 0.00114f
C2710 VPWR.n745 VGND 0.00687f
C2711 VPWR.n746 VGND 0.005442f
C2712 VPWR.n747 VGND 0.020369f
C2713 VPWR.n748 VGND 0.003551f
C2714 VPWR.n749 VGND 0.003278f
C2715 VPWR.n750 VGND 0.003278f
C2716 VPWR.n751 VGND 0.005211f
C2717 VPWR.n752 VGND 0.007102f
C2718 VPWR.n753 VGND 0.007102f
C2719 VPWR.n754 VGND 0.003278f
C2720 VPWR.n755 VGND 0.003278f
C2721 VPWR.n756 VGND 0.003278f
C2722 VPWR.n757 VGND 0.007102f
C2723 VPWR.n758 VGND 0.00687f
C2724 VPWR.t121 VGND 0.003052f
C2725 VPWR.n759 VGND 0.003857f
C2726 VPWR.t256 VGND 0.003062f
C2727 VPWR.n760 VGND 0.004215f
C2728 VPWR.n761 VGND 0.001351f
C2729 VPWR.n762 VGND 0.001942f
C2730 VPWR.n763 VGND 0.001639f
C2731 VPWR.n764 VGND 0.001764f
C2732 VPWR.t313 VGND 0.001373f
C2733 VPWR.t37 VGND 0.001039f
C2734 VPWR.n765 VGND 0.002611f
C2735 VPWR.n766 VGND 0.001247f
C2736 VPWR.t49 VGND 0.003514f
C2737 VPWR.n767 VGND 0.001829f
C2738 VPWR.n768 VGND 0.001099f
C2739 VPWR.n770 VGND 8.79e-19
C2740 VPWR.n771 VGND 8.19e-19
C2741 VPWR.n772 VGND 0.00114f
C2742 VPWR.t531 VGND 0.016311f
C2743 VPWR.t51 VGND 0.001373f
C2744 VPWR.t15 VGND 0.001039f
C2745 VPWR.n773 VGND 0.002435f
C2746 VPWR.n774 VGND 0.002889f
C2747 VPWR.n775 VGND 0.00145f
C2748 VPWR.n776 VGND 0.001139f
C2749 VPWR.t140 VGND 0.002774f
C2750 VPWR.n777 VGND 0.004792f
C2751 VPWR.n778 VGND 0.004583f
C2752 VPWR.n779 VGND 5.17e-19
C2753 VPWR.n780 VGND 0.001099f
C2754 VPWR.n781 VGND 0.00196f
C2755 VPWR.n782 VGND 0.001911f
C2756 VPWR.n783 VGND 0.0017f
C2757 VPWR.n784 VGND 8.22e-19
C2758 VPWR.n785 VGND 0.001942f
C2759 VPWR.t43 VGND 0.003504f
C2760 VPWR.n786 VGND 0.006772f
C2761 VPWR.n787 VGND 0.00145f
C2762 VPWR.t45 VGND 0.001373f
C2763 VPWR.t369 VGND 0.001039f
C2764 VPWR.n788 VGND 0.002435f
C2765 VPWR.t450 VGND 8.5e-19
C2766 VPWR.t47 VGND 8.5e-19
C2767 VPWR.n789 VGND 0.001889f
C2768 VPWR.n790 VGND 0.005112f
C2769 VPWR.t81 VGND 6.39e-19
C2770 VPWR.t481 VGND 1.59e-19
C2771 VPWR.n791 VGND 0.00358f
C2772 VPWR.t18 VGND 6.24e-19
C2773 VPWR.t461 VGND 2.58e-19
C2774 VPWR.n792 VGND 0.003251f
C2775 VPWR.n793 VGND 0.003261f
C2776 VPWR.n794 VGND 0.001942f
C2777 VPWR.t371 VGND 4.21e-19
C2778 VPWR.t424 VGND 4.21e-19
C2779 VPWR.n795 VGND 8.5e-19
C2780 VPWR.n796 VGND 8.8e-19
C2781 VPWR.n797 VGND 2.87e-19
C2782 VPWR.t395 VGND 6.39e-19
C2783 VPWR.t477 VGND 1.59e-19
C2784 VPWR.n798 VGND 0.003565f
C2785 VPWR.n799 VGND 0.003042f
C2786 VPWR.t483 VGND 0.00154f
C2787 VPWR.t195 VGND 0.002774f
C2788 VPWR.n800 VGND 0.004886f
C2789 VPWR.n801 VGND 8.19e-19
C2790 VPWR.n802 VGND 0.00114f
C2791 VPWR.n803 VGND 8.79e-19
C2792 VPWR.n804 VGND 0.001099f
C2793 VPWR.n805 VGND 0.001099f
C2794 VPWR.n806 VGND 0.001716f
C2795 VPWR.n807 VGND 0.001895f
C2796 VPWR.n808 VGND 0.00196f
C2797 VPWR.n809 VGND 0.001461f
C2798 VPWR.t511 VGND 0.016311f
C2799 VPWR.n810 VGND 0.022141f
C2800 VPWR.t237 VGND 0.002797f
C2801 VPWR.t544 VGND 0.005936f
C2802 VPWR.n812 VGND 0.01522f
C2803 VPWR.t238 VGND 0.002797f
C2804 VPWR.n813 VGND 0.007527f
C2805 VPWR.n814 VGND 0.010973f
C2806 VPWR.t196 VGND 0.002774f
C2807 VPWR.n815 VGND 0.004886f
C2808 VPWR.t167 VGND 0.002797f
C2809 VPWR.t517 VGND 0.005936f
C2810 VPWR.n817 VGND 0.01522f
C2811 VPWR.t168 VGND 0.002797f
C2812 VPWR.n818 VGND 0.00829f
C2813 VPWR.t218 VGND 0.002797f
C2814 VPWR.t493 VGND 0.005936f
C2815 VPWR.n820 VGND 0.01522f
C2816 VPWR.t219 VGND 0.002797f
C2817 VPWR.n821 VGND 0.00829f
C2818 VPWR.n822 VGND 0.002757f
C2819 VPWR.n823 VGND 0.006988f
C2820 VPWR.n824 VGND 0.003045f
C2821 VPWR.n825 VGND 0.001942f
C2822 VPWR.n826 VGND 0.003278f
C2823 VPWR.n827 VGND 0.002458f
C2824 VPWR.n828 VGND 0.008604f
C2825 VPWR.n829 VGND 0.008604f
C2826 VPWR.n830 VGND 4.81e-19
C2827 VPWR.n831 VGND 0.001321f
C2828 VPWR.n832 VGND 0.001716f
C2829 VPWR.n833 VGND 0.001895f
C2830 VPWR.n834 VGND 0.00196f
C2831 VPWR.n835 VGND 8.79e-19
C2832 VPWR.n836 VGND 0.001099f
C2833 VPWR.n837 VGND 0.001639f
C2834 VPWR.n838 VGND 0.00114f
C2835 VPWR.n839 VGND 0.003265f
C2836 VPWR.n840 VGND 0.002553f
C2837 VPWR.n841 VGND 2.33e-19
C2838 VPWR.n842 VGND 0.001817f
C2839 VPWR.n843 VGND 0.003278f
C2840 VPWR.n844 VGND 0.002458f
C2841 VPWR.n845 VGND 0.003587f
C2842 VPWR.n846 VGND 0.002972f
C2843 VPWR.n847 VGND 0.001116f
C2844 VPWR.n848 VGND 0.001032f
C2845 VPWR.n849 VGND 0.003278f
C2846 VPWR.n850 VGND 0.003278f
C2847 VPWR.n851 VGND 0.002458f
C2848 VPWR.n852 VGND 4.35e-19
C2849 VPWR.n853 VGND 0.003444f
C2850 VPWR.n854 VGND 5.3e-19
C2851 VPWR.n855 VGND 0.002458f
C2852 VPWR.n856 VGND 0.002458f
C2853 VPWR.n857 VGND 7.44e-19
C2854 VPWR.n858 VGND 0.001829f
C2855 VPWR.n859 VGND 0.002889f
C2856 VPWR.n860 VGND 0.001139f
C2857 VPWR.t141 VGND 0.002774f
C2858 VPWR.n861 VGND 0.004792f
C2859 VPWR.n862 VGND 0.008043f
C2860 VPWR.n863 VGND 0.003278f
C2861 VPWR.n864 VGND 0.002458f
C2862 VPWR.n865 VGND 6.06e-19
C2863 VPWR.n866 VGND 0.008604f
C2864 VPWR.n867 VGND 0.022141f
C2865 VPWR.n868 VGND 0.001639f
C2866 VPWR.n869 VGND 0.001099f
C2867 VPWR.n870 VGND 8.79e-19
C2868 VPWR.n871 VGND 0.00196f
C2869 VPWR.n872 VGND 0.001911f
C2870 VPWR.n873 VGND 0.0017f
C2871 VPWR.n874 VGND 4.3e-19
C2872 VPWR.n875 VGND 9.98e-19
C2873 VPWR.n876 VGND 7.07e-19
C2874 VPWR.n877 VGND 0.003834f
C2875 VPWR.n878 VGND 0.00484f
C2876 VPWR.n879 VGND 0.006486f
C2877 VPWR.t166 VGND 0.028988f
C2878 VPWR.t236 VGND 0.025943f
C2879 VPWR.t194 VGND 0.01754f
C2880 VPWR.t430 VGND 0.021111f
C2881 VPWR.t334 VGND 0.016805f
C2882 VPWR.t476 VGND 0.006722f
C2883 VPWR.t482 VGND 0.010188f
C2884 VPWR.t394 VGND 0.019115f
C2885 VPWR.t423 VGND 0.017855f
C2886 VPWR.t370 VGND 0.012288f
C2887 VPWR.t309 VGND 0.009978f
C2888 VPWR.t17 VGND 0.008823f
C2889 VPWR.t398 VGND 0.009978f
C2890 VPWR.t460 VGND 0.008823f
C2891 VPWR.t480 VGND 0.014389f
C2892 VPWR.t80 VGND 0.015545f
C2893 VPWR.t46 VGND 0.014599f
C2894 VPWR.t449 VGND 0.012499f
C2895 VPWR.t368 VGND 0.009663f
C2896 VPWR.t44 VGND 0.01607f
C2897 VPWR.t42 VGND 0.018695f
C2898 VPWR.t139 VGND 0.013129f
C2899 VPWR.t14 VGND 0.01691f
C2900 VPWR.t50 VGND 0.012604f
C2901 VPWR.t48 VGND 0.009453f
C2902 VPWR.t36 VGND 0.009873f
C2903 VPWR.t312 VGND 0.011238f
C2904 VPWR.n880 VGND 0.010633f
C2905 VPWR.t310 VGND 0.007877f
C2906 VPWR.t254 VGND 0.054931f
C2907 VPWR.t119 VGND 0.061023f
C2908 VPWR.t154 VGND 0.054931f
C2909 VPWR.t174 VGND 0.061023f
C2910 VPWR.n881 VGND 0.027758f
C2911 VPWR.n882 VGND 0.012575f
C2912 VPWR.n883 VGND 7.48e-19
C2913 VPWR.n884 VGND 8.19e-19
C2914 VPWR.n885 VGND 0.001099f
C2915 VPWR.n886 VGND 0.001716f
C2916 VPWR.n887 VGND 0.001895f
C2917 VPWR.n888 VGND 0.129213f
C2918 VPWR.n889 VGND 0.00196f
C2919 VPWR.n890 VGND 0.004028f
C2920 VPWR.n891 VGND 0.001099f
C2921 VPWR.n892 VGND 8.79e-19
C2922 VPWR.t134 VGND 0.041697f
C2923 VPWR.t151 VGND 0.050099f
C2924 VPWR.t163 VGND 0.007877f
C2925 VPWR.t213 VGND 0.054931f
C2926 VPWR.t160 VGND 0.061023f
C2927 VPWR.t110 VGND 0.054931f
C2928 VPWR.t182 VGND 0.061023f
C2929 VPWR.n893 VGND 0.037365f
C2930 VPWR.t239 VGND 0.002797f
C2931 VPWR.t496 VGND 0.005936f
C2932 VPWR.n895 VGND 0.01522f
C2933 VPWR.t240 VGND 0.002797f
C2934 VPWR.n896 VGND 0.00829f
C2935 VPWR.t135 VGND 0.002797f
C2936 VPWR.t519 VGND 0.005936f
C2937 VPWR.n898 VGND 0.01522f
C2938 VPWR.t136 VGND 0.002797f
C2939 VPWR.n899 VGND 0.00829f
C2940 VPWR.n900 VGND 0.00683f
C2941 VPWR.t526 VGND 0.011578f
C2942 VPWR.t152 VGND 0.002804f
C2943 VPWR.n901 VGND 0.016794f
C2944 VPWR.t153 VGND 0.002945f
C2945 VPWR.n902 VGND 0.018712f
C2946 VPWR.n903 VGND 0.00214f
C2947 VPWR.n904 VGND 0.003649f
C2948 VPWR.n905 VGND 0.006048f
C2949 VPWR.n906 VGND 0.007142f
C2950 VPWR.t506 VGND 0.020814f
C2951 VPWR.t164 VGND 0.002774f
C2952 VPWR.n907 VGND 0.034853f
C2953 VPWR.n908 VGND 0.027619f
C2954 VPWR.n909 VGND 0.008727f
C2955 VPWR.n910 VGND 7.48e-19
C2956 VPWR.n911 VGND 8.19e-19
C2957 VPWR.n912 VGND 0.001099f
C2958 VPWR.n913 VGND 0.001716f
C2959 VPWR.n914 VGND 0.001895f
C2960 VPWR.n915 VGND 0.129213f
C2961 VPWR.n916 VGND 0.001895f
C2962 VPWR.n917 VGND 0.001716f
C2963 VPWR.n918 VGND 0.001099f
C2964 VPWR.n919 VGND 0.001461f
C2965 VPWR.n920 VGND 0.00114f
C2966 VPWR.n921 VGND 0.006269f
C2967 VPWR.n922 VGND 0.009053f
C2968 VPWR.t111 VGND 0.003052f
C2969 VPWR.n923 VGND 0.002197f
C2970 VPWR.n924 VGND 0.002586f
C2971 VPWR.n925 VGND 0.002458f
C2972 VPWR.n926 VGND 0.003278f
C2973 VPWR.n927 VGND 0.005211f
C2974 VPWR.n928 VGND 0.007102f
C2975 VPWR.t527 VGND 0.040428f
C2976 VPWR.n929 VGND 0.020369f
C2977 VPWR.n930 VGND 0.005442f
C2978 VPWR.n931 VGND 0.003278f
C2979 VPWR.n932 VGND 0.003278f
C2980 VPWR.n933 VGND 0.003278f
C2981 VPWR.n934 VGND 0.007102f
C2982 VPWR.n935 VGND 0.007102f
C2983 VPWR.n936 VGND 0.00687f
C2984 VPWR.n937 VGND 0.003278f
C2985 VPWR.n938 VGND 0.001942f
C2986 VPWR.n939 VGND 0.00323f
C2987 VPWR.n940 VGND 0.003204f
C2988 VPWR.t161 VGND 0.003052f
C2989 VPWR.n941 VGND 0.003857f
C2990 VPWR.n942 VGND 0.006639f
C2991 VPWR.n943 VGND 0.003278f
C2992 VPWR.n944 VGND 0.001817f
C2993 VPWR.n945 VGND 0.00323f
C2994 VPWR.t214 VGND 0.003052f
C2995 VPWR.n946 VGND 0.002197f
C2996 VPWR.n947 VGND 0.003204f
C2997 VPWR.n948 VGND 0.00114f
C2998 VPWR.n949 VGND 0.001336f
C2999 VPWR.n950 VGND 0.001099f
C3000 VPWR.n951 VGND 0.001716f
C3001 VPWR.n952 VGND 0.001895f
C3002 VPWR.n953 VGND 0.00196f
C3003 VPWR.n954 VGND 0.00196f
C3004 VPWR.n955 VGND 0.001895f
C3005 VPWR.n956 VGND 0.001716f
C3006 VPWR.n957 VGND 0.001099f
C3007 VPWR.n958 VGND 0.001461f
C3008 VPWR.n959 VGND 0.00114f
C3009 VPWR.n960 VGND 0.005211f
C3010 VPWR.n961 VGND 0.007102f
C3011 VPWR.t494 VGND 0.040428f
C3012 VPWR.n962 VGND 0.020369f
C3013 VPWR.n963 VGND 0.005442f
C3014 VPWR.n964 VGND 0.003278f
C3015 VPWR.n965 VGND 0.003278f
C3016 VPWR.n966 VGND 0.003278f
C3017 VPWR.n967 VGND 0.007102f
C3018 VPWR.n968 VGND 0.007102f
C3019 VPWR.n969 VGND 0.00687f
C3020 VPWR.n970 VGND 0.003278f
C3021 VPWR.n971 VGND 0.001942f
C3022 VPWR.n972 VGND 0.00323f
C3023 VPWR.n973 VGND 0.003204f
C3024 VPWR.t158 VGND 0.003052f
C3025 VPWR.n974 VGND 0.003857f
C3026 VPWR.n975 VGND 0.006639f
C3027 VPWR.n976 VGND 0.003278f
C3028 VPWR.n977 VGND 0.001942f
C3029 VPWR.n978 VGND 0.003349f
C3030 VPWR.n979 VGND 0.008563f
C3031 VPWR.n980 VGND 0.001764f
C3032 VPWR.n981 VGND 0.001247f
C3033 VPWR.n982 VGND 0.002837f
C3034 VPWR.n983 VGND 0.004983f
C3035 VPWR.t226 VGND 0.002774f
C3036 VPWR.n984 VGND 0.006371f
C3037 VPWR.n985 VGND 0.025015f
C3038 VPWR.n986 VGND 0.001817f
C3039 VPWR.n987 VGND 0.001321f
C3040 VPWR.n988 VGND 0.001099f
C3041 VPWR.n989 VGND 8.79e-19
C3042 VPWR.n990 VGND 0.00114f
C3043 VPWR.n991 VGND 0.001461f
C3044 VPWR.n992 VGND 0.001099f
C3045 VPWR.n993 VGND 0.001716f
C3046 VPWR.n994 VGND 0.001895f
C3047 VPWR.n995 VGND 0.129213f
C3048 VPWR.n996 VGND 0.001895f
C3049 VPWR.n997 VGND 0.001716f
C3050 VPWR.n998 VGND 0.001099f
C3051 VPWR.n999 VGND 0.001461f
C3052 VPWR.n1000 VGND 0.00114f
C3053 VPWR.n1001 VGND 0.011575f
C3054 VPWR.n1002 VGND 0.011197f
C3055 VPWR.t227 VGND 0.002774f
C3056 VPWR.n1003 VGND 0.006371f
C3057 VPWR.n1004 VGND 0.004216f
C3058 VPWR.n1005 VGND 0.001942f
C3059 VPWR.n1006 VGND 0.001122f
C3060 VPWR.n1007 VGND 9.2e-19
C3061 VPWR.t223 VGND 0.003063f
C3062 VPWR.n1008 VGND 0.003444f
C3063 VPWR.n1009 VGND 0.00348f
C3064 VPWR.n1010 VGND 0.002975f
C3065 VPWR.n1011 VGND 0.003278f
C3066 VPWR.n1012 VGND 0.001942f
C3067 VPWR.n1013 VGND 0.003166f
C3068 VPWR.n1014 VGND 0.018883f
C3069 VPWR.n1015 VGND 0.002896f
C3070 VPWR.n1016 VGND 0.002458f
C3071 VPWR.n1017 VGND 0.003278f
C3072 VPWR.n1018 VGND 0.0022f
C3073 VPWR.n1019 VGND 0.004131f
C3074 VPWR.n1020 VGND 0.003435f
C3075 VPWR.n1021 VGND 0.003278f
C3076 VPWR.n1022 VGND 0.001942f
C3077 VPWR.n1023 VGND 0.002762f
C3078 VPWR.n1024 VGND 0.004131f
C3079 VPWR.t479 VGND 6.39e-19
C3080 VPWR.t308 VGND 1.59e-19
C3081 VPWR.n1025 VGND 0.003565f
C3082 VPWR.n1026 VGND 0.004393f
C3083 VPWR.n1027 VGND 0.003368f
C3084 VPWR.n1028 VGND 0.003278f
C3085 VPWR.n1029 VGND 0.001817f
C3086 VPWR.n1030 VGND 0.001714f
C3087 VPWR.n1031 VGND 0.00114f
C3088 VPWR.t83 VGND 0.001039f
C3089 VPWR.t410 VGND 0.00141f
C3090 VPWR.n1032 VGND 0.002645f
C3091 VPWR.t146 VGND 0.002797f
C3092 VPWR.t528 VGND 0.005936f
C3093 VPWR.n1034 VGND 0.01522f
C3094 VPWR.t147 VGND 0.002797f
C3095 VPWR.n1035 VGND 0.00829f
C3096 VPWR.t408 VGND 0.004348f
C3097 VPWR.t404 VGND 0.001039f
C3098 VPWR.t406 VGND 0.001039f
C3099 VPWR.n1036 VGND 0.002108f
C3100 VPWR.n1037 VGND 0.006261f
C3101 VPWR.n1038 VGND 0.004788f
C3102 VPWR.n1039 VGND 0.001461f
C3103 VPWR.n1040 VGND 0.001336f
C3104 VPWR.n1041 VGND 0.001099f
C3105 VPWR.n1042 VGND 0.00196f
C3106 VPWR.n1043 VGND 8.79e-19
C3107 VPWR.n1044 VGND 0.001099f
C3108 VPWR.n1045 VGND 0.001716f
C3109 VPWR.n1046 VGND 0.001321f
C3110 VPWR.t123 VGND 0.002797f
C3111 VPWR.t535 VGND 0.005936f
C3112 VPWR.n1048 VGND 0.01522f
C3113 VPWR.t124 VGND 0.002797f
C3114 VPWR.n1049 VGND 0.00829f
C3115 VPWR.t172 VGND 0.002797f
C3116 VPWR.t503 VGND 0.005936f
C3117 VPWR.n1051 VGND 0.01522f
C3118 VPWR.t173 VGND 0.002797f
C3119 VPWR.n1052 VGND 0.00829f
C3120 VPWR.n1053 VGND 0.006826f
C3121 VPWR.n1054 VGND 0.002757f
C3122 VPWR.n1055 VGND 0.00276f
C3123 VPWR.n1056 VGND 4.81e-19
C3124 VPWR.n1057 VGND 7.44e-19
C3125 VPWR.n1058 VGND 0.005038f
C3126 VPWR.n1059 VGND 9.4e-19
C3127 VPWR.n1060 VGND 6.24e-19
C3128 VPWR.n1061 VGND 0.001336f
C3129 VPWR.n1062 VGND 0.001099f
C3130 VPWR.n1063 VGND 0.001716f
C3131 VPWR.n1064 VGND 0.001895f
C3132 VPWR.n1065 VGND 0.129213f
C3133 VPWR.n1066 VGND 0.00196f
C3134 VPWR.n1067 VGND 8.79e-19
C3135 VPWR.n1068 VGND 0.001099f
C3136 VPWR.n1069 VGND 8.79e-19
C3137 VPWR.n1070 VGND 8.19e-19
C3138 VPWR.n1071 VGND 0.001099f
C3139 VPWR.n1072 VGND 0.001716f
C3140 VPWR.n1073 VGND 0.001895f
C3141 VPWR.n1074 VGND 0.129213f
C3142 VPWR.n1075 VGND 0.001895f
C3143 VPWR.n1076 VGND 0.001716f
C3144 VPWR.n1077 VGND 0.001321f
C3145 VPWR.n1078 VGND 0.002458f
C3146 VPWR.t25 VGND 6.55e-19
C3147 VPWR.t444 VGND 9.65e-19
C3148 VPWR.n1079 VGND 0.002962f
C3149 VPWR.t416 VGND 0.004392f
C3150 VPWR.t228 VGND 0.002797f
C3151 VPWR.t498 VGND 0.005936f
C3152 VPWR.n1081 VGND 0.01522f
C3153 VPWR.t229 VGND 0.002797f
C3154 VPWR.n1082 VGND 0.00829f
C3155 VPWR.t129 VGND 0.002797f
C3156 VPWR.t520 VGND 0.005936f
C3157 VPWR.n1084 VGND 0.01522f
C3158 VPWR.t130 VGND 0.002797f
C3159 VPWR.n1085 VGND 0.00829f
C3160 VPWR.n1086 VGND 0.002757f
C3161 VPWR.n1087 VGND 0.006895f
C3162 VPWR.n1088 VGND 0.004935f
C3163 VPWR.n1089 VGND 0.004262f
C3164 VPWR.n1090 VGND 0.003278f
C3165 VPWR.n1091 VGND 0.003278f
C3166 VPWR.n1092 VGND 0.001817f
C3167 VPWR.n1093 VGND 7.57e-19
C3168 VPWR.n1094 VGND 0.004855f
C3169 VPWR.n1095 VGND 0.00564f
C3170 VPWR.n1096 VGND 0.001016f
C3171 VPWR.n1097 VGND 0.001817f
C3172 VPWR.n1098 VGND 0.002458f
C3173 VPWR.n1099 VGND 0.002458f
C3174 VPWR.n1100 VGND 0.001009f
C3175 VPWR.n1101 VGND 0.00306f
C3176 VPWR.n1102 VGND 0.00452f
C3177 VPWR.n1103 VGND 0.0119f
C3178 VPWR.n1104 VGND 8.33e-19
C3179 VPWR.n1105 VGND 0.002957f
C3180 VPWR.n1106 VGND 0.00114f
C3181 VPWR.n1107 VGND 0.002458f
C3182 VPWR.n1108 VGND 8.27e-19
C3183 VPWR.n1109 VGND 0.00306f
C3184 VPWR.n1110 VGND 0.004524f
C3185 VPWR.n1111 VGND 9.39e-19
C3186 VPWR.n1112 VGND 0.002458f
C3187 VPWR.n1113 VGND 6.06e-19
C3188 VPWR.n1114 VGND 0.003379f
C3189 VPWR.n1115 VGND 0.005636f
C3190 VPWR.n1116 VGND 0.003359f
C3191 VPWR.n1117 VGND 0.003045f
C3192 VPWR.t118 VGND 0.002797f
C3193 VPWR.n1118 VGND 0.004863f
C3194 VPWR.n1119 VGND 0.007248f
C3195 VPWR.n1120 VGND 0.003278f
C3196 VPWR.n1121 VGND 0.002458f
C3197 VPWR.n1122 VGND 0.003258f
C3198 VPWR.n1123 VGND 0.003685f
C3199 VPWR.n1124 VGND 0.006119f
C3200 VPWR.n1125 VGND 0.001247f
C3201 VPWR.n1126 VGND 0.001122f
C3202 VPWR.n1127 VGND 0.001942f
C3203 VPWR.n1128 VGND 0.003288f
C3204 VPWR.t181 VGND 0.002774f
C3205 VPWR.n1129 VGND 0.00194f
C3206 VPWR.n1130 VGND 0.007844f
C3207 VPWR.n1131 VGND 0.007248f
C3208 VPWR.n1132 VGND 0.005799f
C3209 VPWR.n1133 VGND 0.003278f
C3210 VPWR.n1134 VGND 0.002458f
C3211 VPWR.n1135 VGND 0.001247f
C3212 VPWR.n1136 VGND 0.001018f
C3213 VPWR.n1137 VGND 0.001714f
C3214 VPWR.n1138 VGND 0.001942f
C3215 VPWR.n1139 VGND 0.003278f
C3216 VPWR.n1140 VGND 0.002582f
C3217 VPWR.n1141 VGND 0.005888f
C3218 VPWR.n1142 VGND 0.00348f
C3219 VPWR.n1143 VGND 0.002784f
C3220 VPWR.n1144 VGND 0.001817f
C3221 VPWR.n1145 VGND 0.001321f
C3222 VPWR.n1146 VGND 0.001099f
C3223 VPWR.n1147 VGND 0.00196f
C3224 VPWR.n1148 VGND 8.79e-19
C3225 VPWR.n1149 VGND 0.001716f
C3226 VPWR.n1150 VGND 0.001099f
C3227 VPWR.n1151 VGND 0.001461f
C3228 VPWR.n1152 VGND 0.00114f
C3229 VPWR.n1153 VGND 0.003413f
C3230 VPWR.n1154 VGND 0.004131f
C3231 VPWR.n1155 VGND 0.00114f
C3232 VPWR.n1156 VGND 8.19e-19
C3233 VPWR.n1157 VGND 0.001099f
C3234 VPWR.n1158 VGND 0.001716f
C3235 VPWR.n1159 VGND 0.001895f
C3236 VPWR.n1160 VGND 0.129213f
C3237 VPWR.n1161 VGND 0.105698f
C3238 VPWR.n1162 VGND 0.001895f
C3239 VPWR.n1163 VGND 0.001716f
C3240 VPWR.n1164 VGND 3.05e-19
C3241 VPWR.n1165 VGND 0.001514f
C3242 VPWR.n1166 VGND 0.002945f
C3243 VPWR.n1167 VGND 0.001528f
C3244 VPWR.n1168 VGND 0.001942f
C3245 VPWR.n1169 VGND 0.002458f
C3246 VPWR.n1170 VGND 0.001942f
C3247 VPWR.n1171 VGND 0.004131f
C3248 VPWR.n1172 VGND 0.0022f
C3249 VPWR.n1173 VGND 0.005594f
C3250 VPWR.n1174 VGND 0.003952f
C3251 VPWR.n1175 VGND 0.003278f
C3252 VPWR.n1176 VGND 0.003278f
C3253 VPWR.n1177 VGND 0.002111f
C3254 VPWR.n1178 VGND 0.003884f
C3255 VPWR.n1179 VGND 0.005851f
C3256 VPWR.n1180 VGND 0.001212f
C3257 VPWR.n1181 VGND 0.002458f
C3258 VPWR.n1182 VGND 0.001942f
C3259 VPWR.n1183 VGND 0.003166f
C3260 VPWR.n1184 VGND 0.0022f
C3261 VPWR.n1185 VGND 0.005594f
C3262 VPWR.n1186 VGND 0.003862f
C3263 VPWR.n1187 VGND 0.003278f
C3264 VPWR.n1188 VGND 0.002458f
C3265 VPWR.n1189 VGND 0.001593f
C3266 VPWR.n1190 VGND 8.51e-19
C3267 VPWR.n1191 VGND 6.06e-19
C3268 VPWR.n1192 VGND 8.22e-19
C3269 VPWR.n1193 VGND 0.001716f
C3270 VPWR.n1194 VGND 0.001895f
C3271 VPWR.n1195 VGND 0.00196f
C3272 VPWR.n1196 VGND 8.79e-19
C3273 VPWR.n1197 VGND 0.001099f
.ends

