magic
tech sky130A
magscale 1 2
timestamp 1750693945
<< viali >>
rect 2270 94 2366 128
rect 1340 -694 1458 -658
rect 3116 -702 3248 -664
rect 1288 -2214 1450 -2180
rect 3068 -2212 3214 -2178
rect 2168 -3238 2330 -3200
<< metal1 >>
rect 1672 546 1678 762
rect 1894 546 2412 762
rect 2196 436 2412 546
rect 1378 342 3216 436
rect 1378 262 3218 342
rect 1378 -638 1451 262
rect 2286 160 2359 262
rect 2625 232 2698 262
rect 2260 128 2380 160
rect 2619 159 2625 232
rect 2698 159 2704 232
rect 2260 94 2270 128
rect 2366 94 2380 128
rect 2260 78 2380 94
rect 2086 -12 2374 48
rect 2086 -108 2146 -12
rect 1750 -168 1756 -108
rect 1816 -168 2146 -108
rect 2328 -118 2338 -48
rect 2410 -118 2420 -48
rect 2086 -274 2146 -168
rect 2218 -244 2228 -164
rect 2300 -188 2310 -164
rect 2234 -246 2244 -244
rect 2304 -246 2314 -188
rect 2086 -334 2368 -274
rect 2086 -336 2146 -334
rect 1326 -658 1472 -638
rect 3145 -640 3218 262
rect 1326 -694 1340 -658
rect 1458 -694 1472 -658
rect 1326 -706 1472 -694
rect 3102 -664 3264 -640
rect 3102 -702 3116 -664
rect 3248 -702 3264 -664
rect 3102 -708 3264 -702
rect 923 -736 983 -734
rect 2728 -736 2795 -731
rect 923 -801 1482 -736
rect 923 -803 1481 -801
rect 2728 -803 3280 -736
rect 923 -1064 983 -803
rect 1252 -916 1262 -832
rect 1326 -838 1336 -832
rect 1328 -896 1338 -838
rect 1326 -916 1336 -896
rect 1452 -918 1462 -832
rect 1534 -918 1544 -832
rect 1358 -1034 1368 -964
rect 1434 -1034 1444 -964
rect 1362 -1036 1372 -1034
rect 1430 -1036 1440 -1034
rect 923 -1068 1419 -1064
rect 923 -1126 1420 -1068
rect 2728 -1075 2795 -803
rect 3036 -912 3046 -840
rect 3118 -912 3128 -840
rect 3048 -922 3058 -912
rect 3110 -922 3120 -912
rect 3236 -920 3246 -842
rect 3332 -920 3342 -842
rect 3140 -1036 3150 -970
rect 3214 -988 3224 -970
rect 3152 -1040 3162 -1036
rect 3218 -1040 3228 -988
rect 923 -1129 1419 -1126
rect 923 -1740 983 -1129
rect 2728 -1141 3221 -1075
rect 2728 -1333 2795 -1141
rect 2193 -1400 2199 -1333
rect 2266 -1400 2795 -1333
rect 2728 -1721 2795 -1400
rect 923 -1800 1654 -1740
rect 2728 -1788 3425 -1721
rect 923 -1852 983 -1800
rect 576 -1912 983 -1852
rect 1080 -1908 1090 -1830
rect 1156 -1836 1166 -1830
rect 1164 -1892 1174 -1836
rect 1342 -1840 1352 -1830
rect 1416 -1840 1426 -1830
rect 1156 -1908 1166 -1892
rect 1340 -1898 1350 -1840
rect 1420 -1898 1430 -1840
rect 1342 -1910 1352 -1898
rect 1416 -1910 1426 -1898
rect 1594 -1912 1604 -1834
rect 1682 -1912 1692 -1834
rect 923 -2070 983 -1912
rect 1472 -1962 1482 -1956
rect 1536 -1962 1546 -1956
rect 1204 -2036 1214 -1962
rect 1292 -2036 1302 -1962
rect 1462 -2038 1472 -1962
rect 1548 -2038 1558 -1962
rect 2728 -2063 2795 -1788
rect 2872 -1840 2882 -1826
rect 2870 -1902 2880 -1840
rect 2948 -1888 2958 -1826
rect 3126 -1888 3136 -1828
rect 3206 -1888 3216 -1828
rect 3384 -1840 3394 -1826
rect 2938 -1902 2948 -1888
rect 3128 -1900 3138 -1888
rect 3194 -1900 3204 -1888
rect 3382 -1902 3392 -1840
rect 3458 -1886 3468 -1826
rect 3456 -1902 3466 -1886
rect 3002 -1956 3012 -1946
rect 3072 -1956 3082 -1946
rect 3256 -1954 3266 -1950
rect 3328 -1954 3338 -1950
rect 2998 -2032 3008 -1956
rect 3078 -2032 3088 -1956
rect 3246 -2032 3256 -1954
rect 3254 -2034 3264 -2032
rect 3332 -2034 3342 -1954
rect 923 -2130 1634 -2070
rect 2728 -2130 3425 -2063
rect 1525 -2132 1590 -2130
rect 2728 -2131 2795 -2130
rect 1254 -2180 1470 -2170
rect 1254 -2214 1288 -2180
rect 1450 -2214 1470 -2180
rect 1254 -2286 1470 -2214
rect 3056 -2178 3242 -2162
rect 3056 -2212 3068 -2178
rect 3214 -2212 3242 -2178
rect 1291 -3416 1377 -2286
rect 3056 -2292 3242 -2212
rect 1793 -2818 2530 -2756
rect 1793 -2931 1855 -2818
rect 1964 -2926 1974 -2854
rect 2042 -2926 2052 -2854
rect 2234 -2864 2244 -2858
rect 2296 -2864 2306 -2858
rect 2492 -2860 2502 -2856
rect 2558 -2860 2568 -2856
rect 2224 -2928 2234 -2864
rect 2306 -2928 2316 -2864
rect 2482 -2928 2492 -2860
rect 2562 -2928 2572 -2860
rect 1557 -2993 1563 -2931
rect 1625 -2993 1855 -2931
rect 2104 -2988 2114 -2976
rect 2172 -2988 2182 -2976
rect 2360 -2986 2370 -2976
rect 2426 -2986 2436 -2976
rect 1793 -3099 1855 -2993
rect 2100 -3058 2110 -2988
rect 2178 -3058 2188 -2988
rect 2358 -3054 2368 -2986
rect 2436 -3054 2446 -2986
rect 1793 -3161 2503 -3099
rect 2152 -3200 2342 -3190
rect 2152 -3238 2168 -3200
rect 2330 -3238 2342 -3200
rect 2152 -3300 2342 -3238
rect 2223 -3416 2309 -3300
rect 2727 -3359 2733 -3273
rect 2819 -3359 2825 -3273
rect 2733 -3416 2819 -3359
rect 3137 -3416 3223 -2292
rect 1291 -3511 3224 -3416
rect 1292 -3610 3224 -3511
rect 2148 -3754 2348 -3610
rect 2148 -3960 2348 -3954
<< via1 >>
rect 1678 546 1894 762
rect 2625 159 2698 232
rect 1756 -168 1816 -108
rect 2338 -118 2410 -48
rect 2228 -188 2300 -164
rect 2228 -244 2304 -188
rect 2244 -246 2304 -244
rect 1262 -838 1326 -832
rect 1262 -896 1328 -838
rect 1262 -916 1326 -896
rect 1462 -918 1534 -832
rect 1368 -1034 1434 -964
rect 1372 -1036 1430 -1034
rect 3046 -912 3118 -840
rect 3058 -922 3110 -912
rect 3246 -920 3332 -842
rect 3150 -988 3214 -970
rect 3150 -1036 3218 -988
rect 3162 -1040 3218 -1036
rect 2199 -1400 2266 -1333
rect 1090 -1836 1156 -1830
rect 1090 -1892 1164 -1836
rect 1352 -1840 1416 -1830
rect 1090 -1908 1156 -1892
rect 1350 -1898 1420 -1840
rect 1352 -1910 1416 -1898
rect 1604 -1912 1682 -1834
rect 1482 -1962 1536 -1956
rect 1214 -2036 1292 -1962
rect 1472 -2038 1548 -1962
rect 2882 -1840 2948 -1826
rect 2880 -1888 2948 -1840
rect 3136 -1888 3206 -1828
rect 3394 -1840 3458 -1826
rect 2880 -1902 2938 -1888
rect 3138 -1900 3194 -1888
rect 3392 -1886 3458 -1840
rect 3392 -1902 3456 -1886
rect 3012 -1956 3072 -1946
rect 3266 -1954 3328 -1950
rect 3008 -2032 3078 -1956
rect 3256 -2032 3332 -1954
rect 3264 -2034 3332 -2032
rect 1974 -2926 2042 -2854
rect 2244 -2864 2296 -2858
rect 2502 -2860 2558 -2856
rect 2234 -2928 2306 -2864
rect 2492 -2928 2562 -2860
rect 1563 -2993 1625 -2931
rect 2114 -2988 2172 -2976
rect 2370 -2986 2426 -2976
rect 2110 -3058 2178 -2988
rect 2368 -3054 2436 -2986
rect 2733 -3359 2819 -3273
rect 2148 -3954 2348 -3754
<< metal2 >>
rect 1128 763 1337 772
rect 1678 763 1894 768
rect 1337 762 1894 763
rect 1337 554 1678 762
rect 1128 545 1337 554
rect 1518 546 1678 554
rect 1678 540 1894 546
rect 2625 232 2698 238
rect 2625 -34 2698 159
rect 2204 -48 2698 -34
rect 1756 -108 1816 -102
rect 606 -168 1756 -108
rect 2204 -118 2338 -48
rect 2410 -118 2698 -48
rect 2204 -124 2698 -118
rect 2338 -128 2410 -124
rect 1756 -174 1816 -168
rect 2228 -164 2300 -154
rect 2200 -244 2228 -172
rect 2300 -188 2632 -172
rect 2200 -246 2244 -244
rect 2304 -246 2632 -188
rect 2200 -260 2632 -246
rect 1262 -826 1326 -822
rect 1462 -826 1534 -822
rect 2540 -826 2628 -260
rect 1228 -832 2629 -826
rect 1228 -910 1262 -832
rect 1326 -838 1462 -832
rect 1328 -896 1462 -838
rect 1236 -916 1262 -910
rect 1326 -916 1462 -896
rect 1236 -918 1462 -916
rect 1534 -835 2629 -832
rect 3046 -835 3118 -830
rect 3246 -835 3332 -832
rect 1534 -836 3462 -835
rect 1534 -840 3466 -836
rect 1534 -912 3046 -840
rect 3118 -842 3466 -840
rect 3118 -912 3246 -842
rect 1534 -918 3058 -912
rect 1236 -922 3058 -918
rect 3110 -920 3246 -912
rect 3332 -920 3466 -842
rect 3110 -922 3466 -920
rect 1236 -924 3466 -922
rect 1262 -926 1326 -924
rect 1462 -928 1534 -924
rect 3058 -932 3110 -924
rect 3246 -930 3332 -924
rect 1368 -956 1434 -954
rect 1234 -964 1854 -956
rect 3150 -962 3214 -960
rect 1234 -966 1368 -964
rect 1232 -1034 1368 -966
rect 1434 -976 1854 -964
rect 1434 -1034 1771 -976
rect 1232 -1036 1372 -1034
rect 1430 -1036 1771 -1034
rect 1232 -1049 1771 -1036
rect 1844 -1048 1854 -976
rect 3058 -970 3798 -962
rect 3058 -1036 3150 -970
rect 3214 -972 3798 -970
rect 3214 -988 3800 -972
rect 3058 -1040 3162 -1036
rect 3218 -1040 3800 -988
rect 3058 -1045 3800 -1040
rect 3058 -1048 3798 -1045
rect 1844 -1049 1853 -1048
rect 1232 -1056 1852 -1049
rect 3162 -1050 3218 -1048
rect 2199 -1333 2266 -1327
rect 559 -1400 2199 -1333
rect 2199 -1406 2266 -1400
rect 1090 -1828 1156 -1820
rect 1352 -1828 1416 -1820
rect 1604 -1828 1682 -1824
rect 2834 -1826 3829 -1820
rect 1064 -1830 1868 -1828
rect 1064 -1908 1090 -1830
rect 1156 -1836 1352 -1830
rect 1164 -1840 1352 -1836
rect 1416 -1834 1868 -1830
rect 1416 -1840 1604 -1834
rect 1164 -1892 1350 -1840
rect 1156 -1898 1350 -1892
rect 1420 -1898 1604 -1840
rect 1156 -1908 1352 -1898
rect 1064 -1910 1352 -1908
rect 1416 -1910 1604 -1898
rect 1064 -1912 1604 -1910
rect 1682 -1912 1868 -1834
rect 1952 -1912 1961 -1828
rect 2834 -1840 2882 -1826
rect 2948 -1828 3394 -1826
rect 2834 -1902 2880 -1840
rect 2948 -1888 3136 -1828
rect 3206 -1840 3394 -1828
rect 3458 -1836 3829 -1826
rect 3206 -1888 3392 -1840
rect 3458 -1886 3830 -1836
rect 2938 -1900 3138 -1888
rect 3194 -1900 3392 -1888
rect 2938 -1902 3392 -1900
rect 3456 -1902 3830 -1886
rect 2834 -1908 3830 -1902
rect 2880 -1912 2938 -1908
rect 3138 -1910 3194 -1908
rect 3392 -1912 3456 -1908
rect 1090 -1918 1156 -1912
rect 1352 -1920 1416 -1912
rect 1604 -1922 1682 -1912
rect 3012 -1946 3072 -1936
rect 3266 -1944 3328 -1940
rect 1482 -1950 1536 -1946
rect 3008 -1950 3012 -1946
rect 1070 -1956 3012 -1950
rect 3072 -1950 3078 -1946
rect 3256 -1950 3332 -1944
rect 3072 -1954 3266 -1950
rect 3328 -1954 3604 -1950
rect 3072 -1956 3256 -1954
rect 1066 -1962 1482 -1956
rect 1536 -1962 3008 -1956
rect 1066 -2036 1214 -1962
rect 1292 -2036 1472 -1962
rect 1066 -2038 1472 -2036
rect 1548 -2032 3008 -1962
rect 3078 -2032 3256 -1956
rect 1548 -2034 3264 -2032
rect 3332 -2034 3604 -1954
rect 1548 -2036 3604 -2034
rect 1548 -2038 2414 -2036
rect 1066 -2054 2414 -2038
rect 3008 -2042 3078 -2036
rect 3256 -2042 3332 -2036
rect 3264 -2044 3332 -2042
rect 1068 -2056 2414 -2054
rect 1974 -2846 2042 -2844
rect 2290 -2846 2414 -2056
rect 1932 -2854 2626 -2846
rect 1563 -2931 1625 -2925
rect 667 -2993 1563 -2931
rect 1932 -2926 1974 -2854
rect 2042 -2856 2626 -2854
rect 2042 -2858 2502 -2856
rect 2042 -2864 2244 -2858
rect 2296 -2860 2502 -2858
rect 2558 -2860 2626 -2856
rect 2296 -2864 2492 -2860
rect 2042 -2926 2234 -2864
rect 1932 -2928 2234 -2926
rect 2306 -2928 2492 -2864
rect 2562 -2928 2626 -2860
rect 1932 -2934 2626 -2928
rect 1974 -2936 2042 -2934
rect 2234 -2938 2306 -2934
rect 2492 -2938 2562 -2934
rect 1563 -2999 1625 -2993
rect 2050 -2976 2818 -2966
rect 2050 -2988 2114 -2976
rect 2172 -2986 2370 -2976
rect 2426 -2980 2818 -2976
rect 2426 -2986 2819 -2980
rect 2172 -2988 2368 -2986
rect 2050 -3058 2110 -2988
rect 2178 -3054 2368 -2988
rect 2436 -3054 2819 -2986
rect 2178 -3058 2819 -3054
rect 2050 -3066 2819 -3058
rect 2110 -3068 2178 -3066
rect 2733 -3273 2819 -3066
rect 2733 -3365 2819 -3359
rect 1788 -3965 1797 -3751
rect 2011 -3754 2192 -3751
rect 2011 -3954 2148 -3754
rect 2348 -3954 2354 -3754
rect 2011 -3965 2192 -3954
<< via2 >>
rect 1128 554 1337 763
rect 1771 -1049 1844 -976
rect 1868 -1912 1952 -1828
rect 1797 -3965 2011 -3751
<< metal3 >>
rect 1123 763 1342 768
rect 1123 554 1128 763
rect 1337 554 1342 763
rect 1123 549 1342 554
rect 1128 523 1337 549
rect 1128 308 1337 314
rect 1771 -521 3804 -448
rect 1771 -971 1844 -521
rect 1766 -976 1849 -971
rect 1766 -1049 1771 -976
rect 1844 -1049 1849 -976
rect 1766 -1054 1849 -1049
rect 1863 -1828 1957 -1823
rect 1863 -1912 1868 -1828
rect 1952 -1912 1957 -1828
rect 1863 -1917 1957 -1912
rect 1868 -2294 1952 -1917
rect 1868 -2378 3830 -2294
rect 1792 -3751 2016 -3746
rect 501 -3965 507 -3751
rect 721 -3965 1797 -3751
rect 2011 -3965 2016 -3751
rect 1792 -3970 2016 -3965
<< via3 >>
rect 1128 314 1337 523
rect 507 -3965 721 -3751
<< metal4 >>
rect 516 -3585 716 1564
rect 1127 523 1338 524
rect 1127 314 1128 523
rect 1337 314 1338 523
rect 1127 313 1338 314
rect 507 -3750 721 -3585
rect 506 -3751 722 -3750
rect 506 -3965 507 -3751
rect 721 -3965 722 -3751
rect 506 -3966 722 -3965
rect 1128 -4682 1337 313
use sky130_fd_pr__nfet_01v8_lvt_648S5X  sky130_fd_pr__nfet_01v8_lvt_648S5X_0
timestamp 1749574077
transform 1 0 2321 0 1 -146
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QBKD3  sky130_fd_pr__pfet_01v8_lvt_4QBKD3_1
timestamp 1749574077
transform 1 0 2269 0 1 -2951
box -423 -319 423 319
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  XM1
timestamp 1749574077
transform 1 0 3183 0 1 -940
box -263 -310 263 310
use sky130_fd_pr__pfet_01v8_lvt_4QBKD3  XM10
timestamp 1749574077
transform 1 0 1383 0 1 -1931
box -423 -319 423 319
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  XM11
timestamp 1749574077
transform 1 0 1401 0 1 -932
box -263 -310 263 310
use sky130_fd_pr__pfet_01v8_lvt_4QBKD3  XM12
timestamp 1749574077
transform 1 0 3169 0 1 -1927
box -423 -319 423 319
<< end >>
