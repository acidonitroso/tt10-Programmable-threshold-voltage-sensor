magic
tech sky130A
magscale 1 2
timestamp 1750416658
<< viali >>
rect 552 2158 643 2198
rect 544 960 716 1015
<< metal1 >>
rect 144 2242 668 2318
rect 144 2006 220 2242
rect 531 2198 666 2242
rect 531 2158 552 2198
rect 643 2158 666 2198
rect 531 2150 666 2158
rect 533 2148 664 2150
rect 265 2109 344 2111
rect 144 1924 220 1930
rect 260 2048 742 2109
rect 260 1772 344 2048
rect 448 1999 458 2000
rect 444 1938 454 1999
rect 448 1934 458 1938
rect 518 1934 528 2000
rect 708 1928 718 2000
rect 776 1989 786 2000
rect 711 1927 721 1928
rect 784 1927 794 1989
rect 578 1876 588 1886
rect 652 1876 662 1886
rect 576 1805 586 1876
rect 653 1805 663 1876
rect 260 1711 740 1772
rect 260 1466 344 1711
rect 260 1379 679 1466
rect 260 1117 344 1379
rect 538 1212 548 1288
rect 608 1279 618 1288
rect 609 1223 619 1279
rect 608 1212 618 1223
rect 648 1212 658 1288
rect 716 1234 726 1288
rect 714 1212 724 1234
rect 260 1056 664 1117
rect 530 1015 723 1027
rect 530 960 544 1015
rect 716 960 723 1015
rect 530 942 723 960
rect 402 873 408 941
rect 476 873 482 941
rect 408 783 476 873
rect 563 783 656 942
rect 408 715 656 783
rect 563 698 656 715
<< via1 >>
rect 144 1930 220 2006
rect 458 1999 518 2000
rect 454 1938 518 1999
rect 458 1934 518 1938
rect 718 1989 776 2000
rect 718 1928 784 1989
rect 721 1927 784 1928
rect 588 1876 652 1886
rect 586 1805 653 1876
rect 548 1279 608 1288
rect 548 1223 609 1279
rect 548 1212 608 1223
rect 658 1234 716 1288
rect 658 1212 714 1234
rect 408 873 476 941
<< metal2 >>
rect 458 2009 518 2010
rect 454 2006 518 2009
rect 718 2006 776 2010
rect 138 1930 144 2006
rect 220 2002 790 2006
rect 220 2000 820 2002
rect 220 1999 458 2000
rect 220 1938 454 1999
rect 220 1934 458 1938
rect 518 1934 718 2000
rect 776 1989 820 2000
rect 220 1930 718 1934
rect 138 1928 718 1930
rect 138 1927 721 1928
rect 784 1927 820 1989
rect 138 1924 820 1927
rect 718 1918 784 1924
rect 721 1917 784 1918
rect 588 1890 652 1896
rect 440 1886 672 1890
rect 440 1876 588 1886
rect 652 1882 672 1886
rect 652 1876 1016 1882
rect 440 1870 586 1876
rect 439 1805 586 1870
rect 653 1806 1016 1876
rect 653 1805 1013 1806
rect 439 1804 1013 1805
rect 586 1795 653 1804
rect 410 1289 608 1300
rect 947 1298 1013 1804
rect 410 1288 609 1289
rect 410 1285 548 1288
rect 408 1212 548 1285
rect 608 1279 609 1288
rect 608 1213 609 1223
rect 654 1288 1014 1298
rect 408 1202 608 1212
rect 654 1212 658 1288
rect 716 1234 1014 1288
rect 714 1212 1014 1234
rect 654 1202 1014 1212
rect 408 941 476 1202
rect 408 867 476 873
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM22 ~/tt10-analog-template-psei-def/mag
timestamp 1749574077
transform 1 0 631 0 1 1250
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM25 ~/tt10-analog-template-psei-def/mag
timestamp 1749567790
transform 1 0 619 0 1 1913
box -295 -319 295 319
<< end >>
