magic
tech sky130A
magscale 1 2
timestamp 1750428065
<< viali >>
rect 1226 -156 1372 -122
rect 2244 -164 2390 -128
rect 1248 -1110 1342 -1074
rect 2278 -1116 2382 -1074
rect 1286 -2462 1354 -2428
rect 2312 -2464 2384 -2428
rect 1280 -3236 1378 -3202
rect 2314 -3246 2396 -3206
<< metal1 >>
rect 899 7 2725 17
rect 899 -58 2727 7
rect 899 -290 974 -58
rect 1214 -122 1380 -58
rect 1214 -156 1226 -122
rect 1372 -156 1380 -122
rect 1214 -170 1380 -156
rect 2234 -128 2402 -58
rect 2234 -164 2244 -128
rect 2390 -164 2402 -128
rect 2234 -178 2402 -164
rect 1158 -272 2438 -208
rect 893 -365 899 -341
rect 1136 -314 1146 -300
rect 893 -371 974 -365
rect 893 -939 968 -371
rect 1130 -376 1140 -314
rect 1216 -368 1226 -300
rect 1140 -386 1150 -376
rect 1212 -386 1222 -368
rect 1392 -374 1402 -304
rect 1482 -374 1492 -304
rect 1396 -384 1406 -374
rect 1470 -384 1480 -374
rect 1272 -510 1282 -432
rect 1344 -510 1354 -432
rect 1772 -542 1848 -272
rect 2650 -308 2727 -58
rect 2158 -384 2168 -312
rect 2244 -384 2254 -312
rect 2418 -382 2428 -314
rect 2502 -382 2512 -314
rect 2646 -376 2656 -308
rect 2724 -314 2734 -308
rect 2727 -376 2734 -314
rect 2288 -508 2298 -430
rect 2376 -508 2386 -430
rect 2290 -514 2300 -508
rect 2368 -514 2378 -508
rect 1158 -608 2471 -542
rect 1624 -676 1709 -608
rect 1624 -732 1638 -676
rect 1694 -732 1709 -676
rect 1624 -734 1709 -732
rect 2650 -928 2727 -376
rect 893 -944 1347 -939
rect 893 -1008 1350 -944
rect 2271 -948 2727 -928
rect 2266 -1003 2727 -948
rect 893 -1014 1348 -1008
rect 1236 -1074 1348 -1014
rect 1236 -1110 1248 -1074
rect 1342 -1110 1348 -1074
rect 1236 -1122 1348 -1110
rect 2266 -1074 2392 -1003
rect 2266 -1116 2278 -1074
rect 2382 -1116 2392 -1074
rect 2266 -1130 2392 -1116
rect 1149 -1225 2475 -1158
rect 1142 -1330 1152 -1254
rect 1216 -1330 1226 -1254
rect 1398 -1334 1408 -1258
rect 1490 -1334 1500 -1258
rect 1272 -1452 1282 -1384
rect 1336 -1406 1346 -1384
rect 1274 -1466 1284 -1452
rect 1342 -1466 1352 -1406
rect 1774 -1496 1848 -1225
rect 2162 -1338 2172 -1270
rect 2246 -1338 2256 -1270
rect 2422 -1336 2432 -1270
rect 2504 -1336 2514 -1270
rect 2292 -1468 2302 -1394
rect 2378 -1468 2388 -1394
rect 1164 -1570 2447 -1496
rect 1907 -1815 1981 -1570
rect 1907 -1895 1981 -1889
rect 1242 -2000 2416 -1982
rect 1240 -2054 2417 -2000
rect 1614 -2088 1686 -2054
rect 1236 -2164 1246 -2098
rect 1302 -2164 1312 -2098
rect 1614 -2166 1686 -2160
rect 1332 -2230 1342 -2212
rect 1328 -2290 1338 -2230
rect 1400 -2290 1410 -2212
rect 1764 -2318 1848 -2054
rect 2354 -2156 2364 -2088
rect 2420 -2094 2430 -2088
rect 2356 -2172 2366 -2156
rect 2432 -2162 2442 -2094
rect 2426 -2172 2436 -2162
rect 2262 -2236 2272 -2214
rect 2258 -2290 2268 -2236
rect 2326 -2276 2336 -2214
rect 2322 -2290 2332 -2276
rect 1218 -2386 2380 -2318
rect 1274 -2428 1368 -2414
rect 1274 -2462 1286 -2428
rect 1354 -2462 1368 -2428
rect 1274 -2514 1368 -2462
rect 2302 -2428 2394 -2416
rect 2302 -2464 2312 -2428
rect 2384 -2464 2394 -2428
rect 2302 -2504 2394 -2464
rect 2313 -2511 2383 -2504
rect 1292 -2528 1356 -2514
rect 2313 -2587 2383 -2581
rect 1292 -2598 1356 -2592
rect 1252 -2778 2398 -2756
rect 1250 -2832 2399 -2778
rect 1342 -2874 1352 -2872
rect 1410 -2874 1420 -2872
rect 1338 -2942 1348 -2874
rect 1412 -2942 1422 -2874
rect 1248 -3004 1258 -2984
rect 1310 -3004 1320 -2984
rect 1244 -3060 1254 -3004
rect 1312 -3060 1322 -3004
rect 1503 -3017 1565 -3011
rect 1503 -3096 1565 -3079
rect 1766 -3096 1848 -2832
rect 2272 -2934 2282 -2874
rect 2340 -2934 2350 -2874
rect 2274 -2942 2284 -2934
rect 2336 -2942 2346 -2934
rect 2366 -3068 2376 -2992
rect 2432 -3068 2442 -2992
rect 897 -3225 903 -3155
rect 973 -3225 979 -3155
rect 1254 -3158 2399 -3096
rect 1264 -3202 1402 -3192
rect 903 -3267 973 -3225
rect 1264 -3236 1280 -3202
rect 1378 -3236 1402 -3202
rect 1264 -3267 1402 -3236
rect 2296 -3206 2428 -3192
rect 2296 -3246 2314 -3206
rect 2396 -3246 2428 -3206
rect 2676 -3225 2682 -3158
rect 2749 -3225 2755 -3158
rect 1766 -3267 1772 -3254
rect 903 -3330 1772 -3267
rect 1848 -3267 1854 -3254
rect 2296 -3267 2428 -3246
rect 2682 -3267 2749 -3225
rect 1848 -3330 2749 -3267
rect 903 -3349 2749 -3330
rect 963 -3350 2693 -3349
<< via1 >>
rect 899 -365 974 -290
rect 1146 -314 1216 -300
rect 1140 -368 1216 -314
rect 1140 -376 1212 -368
rect 1150 -386 1212 -376
rect 1402 -374 1482 -304
rect 1406 -384 1470 -374
rect 1282 -510 1344 -432
rect 2168 -384 2244 -312
rect 2428 -382 2502 -314
rect 2656 -314 2724 -308
rect 2656 -376 2727 -314
rect 2298 -508 2376 -430
rect 2300 -514 2368 -508
rect 1638 -732 1694 -676
rect 1152 -1330 1216 -1254
rect 1408 -1334 1490 -1258
rect 1282 -1406 1336 -1384
rect 1282 -1452 1342 -1406
rect 1284 -1466 1342 -1452
rect 2172 -1338 2246 -1270
rect 2432 -1336 2504 -1270
rect 2302 -1468 2378 -1394
rect 1907 -1889 1981 -1815
rect 1246 -2164 1302 -2098
rect 1614 -2160 1686 -2088
rect 1342 -2230 1400 -2212
rect 1338 -2290 1400 -2230
rect 2364 -2094 2420 -2088
rect 2364 -2156 2432 -2094
rect 2366 -2162 2432 -2156
rect 2366 -2172 2426 -2162
rect 2272 -2236 2326 -2214
rect 2268 -2276 2326 -2236
rect 2268 -2290 2322 -2276
rect 1292 -2592 1356 -2528
rect 2313 -2581 2383 -2511
rect 1352 -2874 1410 -2872
rect 1348 -2942 1412 -2874
rect 1258 -3004 1310 -2984
rect 1254 -3060 1312 -3004
rect 1503 -3079 1565 -3017
rect 2282 -2934 2340 -2874
rect 2284 -2942 2336 -2934
rect 2376 -3068 2432 -2992
rect 903 -3225 973 -3155
rect 2682 -3225 2749 -3158
rect 1772 -3330 1848 -3254
<< metal2 >>
rect 893 -292 899 -290
rect 890 -365 899 -292
rect 974 -292 1031 -290
rect 1146 -292 1216 -290
rect 974 -300 1490 -292
rect 974 -314 1146 -300
rect 1216 -304 1490 -300
rect 974 -365 1140 -314
rect 890 -376 1140 -365
rect 1216 -368 1402 -304
rect 1212 -374 1402 -368
rect 1482 -374 1490 -304
rect 2168 -310 2244 -302
rect 2428 -310 2502 -304
rect 2656 -308 2724 -298
rect 890 -386 1150 -376
rect 1212 -384 1406 -374
rect 1470 -384 1490 -374
rect 2162 -312 2656 -310
rect 2162 -384 2168 -312
rect 2244 -314 2656 -312
rect 2724 -314 2734 -310
rect 2244 -382 2428 -314
rect 2502 -376 2656 -314
rect 2727 -376 2734 -314
rect 2502 -382 2734 -376
rect 2244 -384 2734 -382
rect 1212 -386 1490 -384
rect 890 -390 1490 -386
rect 1150 -396 1212 -390
rect 1406 -394 1470 -390
rect 2168 -394 2244 -384
rect 2428 -392 2502 -384
rect 2656 -386 2724 -384
rect 1282 -432 1344 -422
rect 2298 -428 2376 -420
rect 2168 -430 2736 -428
rect 898 -444 1282 -432
rect 897 -506 1282 -444
rect 897 -1254 959 -506
rect 1344 -444 1472 -432
rect 1344 -506 1474 -444
rect 1282 -520 1344 -510
rect 2168 -508 2298 -430
rect 2376 -442 2736 -430
rect 2376 -508 2739 -442
rect 2168 -514 2300 -508
rect 2368 -514 2739 -508
rect 2168 -516 2739 -514
rect 2170 -520 2739 -516
rect 2300 -524 2368 -520
rect 1622 -670 1693 -665
rect 1622 -676 1694 -670
rect 1622 -732 1638 -676
rect 1152 -1254 1216 -1244
rect 1408 -1254 1490 -1248
rect 896 -1330 1152 -1254
rect 1216 -1258 1490 -1254
rect 1216 -1330 1408 -1258
rect 896 -1334 1408 -1330
rect 1490 -1321 1495 -1259
rect 896 -1340 1490 -1334
rect 1408 -1344 1490 -1340
rect 1282 -1380 1336 -1374
rect 1622 -1380 1694 -732
rect 2661 -1267 2739 -520
rect 2161 -1270 2739 -1267
rect 2161 -1338 2172 -1270
rect 2246 -1336 2432 -1270
rect 2504 -1336 2739 -1270
rect 2246 -1338 2739 -1336
rect 2161 -1345 2739 -1338
rect 2172 -1348 2246 -1345
rect 2432 -1346 2504 -1345
rect 898 -1384 1694 -1380
rect 898 -1452 1282 -1384
rect 1336 -1406 1694 -1384
rect 2302 -1394 2378 -1384
rect 898 -1466 1284 -1452
rect 1342 -1466 1694 -1406
rect 898 -1482 1693 -1466
rect 2164 -1468 2302 -1398
rect 2378 -1403 2738 -1398
rect 2378 -1468 2739 -1403
rect 2164 -1474 2739 -1468
rect 2302 -1478 2378 -1474
rect 898 -2090 972 -1482
rect 1901 -1889 1907 -1815
rect 1981 -1889 1987 -1815
rect 1246 -2090 1302 -2088
rect 898 -2098 1397 -2090
rect 898 -2154 1246 -2098
rect 901 -2161 1246 -2154
rect 1302 -2161 1397 -2098
rect 1608 -2160 1614 -2088
rect 1686 -2160 1692 -2088
rect 1246 -2174 1302 -2164
rect 1342 -2208 1400 -2202
rect 898 -2212 1400 -2208
rect 898 -2230 1342 -2212
rect 898 -2290 1338 -2230
rect 1400 -2290 1418 -2228
rect 899 -2294 1418 -2290
rect 899 -2848 965 -2294
rect 1338 -2300 1400 -2294
rect 1614 -2376 1686 -2160
rect 1907 -2187 1981 -1889
rect 2364 -2084 2420 -2078
rect 2668 -2084 2739 -1474
rect 2242 -2088 2739 -2084
rect 2242 -2156 2364 -2088
rect 2420 -2094 2739 -2088
rect 2242 -2166 2366 -2156
rect 2432 -2157 2739 -2094
rect 2432 -2162 2738 -2157
rect 2244 -2172 2366 -2166
rect 2426 -2172 2738 -2162
rect 2366 -2182 2426 -2172
rect 2272 -2214 2326 -2204
rect 1907 -2270 1981 -2261
rect 2254 -2236 2272 -2218
rect 2326 -2229 2746 -2218
rect 2254 -2290 2268 -2236
rect 2326 -2276 2750 -2229
rect 2322 -2290 2750 -2276
rect 2254 -2300 2750 -2290
rect 2258 -2301 2750 -2300
rect 1614 -2457 1686 -2448
rect 1772 -2528 1848 -2522
rect 2307 -2528 2313 -2511
rect 1286 -2592 1292 -2528
rect 1356 -2581 2313 -2528
rect 2383 -2581 2389 -2511
rect 1356 -2592 2388 -2581
rect 899 -2864 1416 -2848
rect 900 -2872 1416 -2864
rect 900 -2874 1352 -2872
rect 1410 -2874 1416 -2872
rect 900 -2942 1348 -2874
rect 1412 -2942 1416 -2874
rect 1348 -2952 1416 -2942
rect 1258 -2980 1310 -2974
rect 904 -2984 1434 -2980
rect 904 -3003 1258 -2984
rect 903 -3004 1258 -3003
rect 1310 -3004 1434 -2984
rect 903 -3060 1254 -3004
rect 1312 -3060 1434 -3004
rect 903 -3070 1434 -3060
rect 1496 -3017 1573 -3009
rect 903 -3073 1433 -3070
rect 903 -3155 973 -3073
rect 903 -3231 973 -3225
rect 1496 -3079 1503 -3017
rect 1565 -3079 1573 -3017
rect 1496 -3500 1573 -3079
rect 1772 -3254 1848 -2592
rect 2678 -2849 2750 -2301
rect 2267 -2850 2751 -2849
rect 2248 -2874 2752 -2850
rect 2248 -2934 2282 -2874
rect 2340 -2934 2752 -2874
rect 2248 -2942 2284 -2934
rect 2336 -2942 2752 -2934
rect 2248 -2946 2752 -2942
rect 2284 -2952 2336 -2946
rect 2376 -2988 2432 -2982
rect 2246 -2992 2750 -2988
rect 2246 -3011 2376 -2992
rect 2245 -3068 2376 -3011
rect 2432 -3068 2750 -2992
rect 2245 -3078 2750 -3068
rect 2246 -3084 2750 -3078
rect 2682 -3158 2749 -3084
rect 2682 -3231 2749 -3225
rect 1772 -3336 1848 -3330
<< via2 >>
rect 1907 -2261 1981 -2187
rect 1614 -2448 1686 -2376
<< metal3 >>
rect 1902 -2187 1986 -2182
rect 1902 -2261 1907 -2187
rect 1981 -2261 1986 -2187
rect 1902 -2266 1986 -2261
rect 1609 -2376 1691 -2371
rect 1609 -2448 1614 -2376
rect 1686 -2448 1691 -2376
rect 1609 -2453 1691 -2448
rect 1614 -3500 1686 -2453
rect 1907 -3499 1981 -2266
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM1
timestamp 1749567790
transform -1 0 1323 0 1 -1361
box -295 -319 295 319
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM2
timestamp 1749567790
transform 1 0 2343 0 1 -413
box -295 -319 295 319
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM3
timestamp 1749567790
transform 1 0 1321 0 1 -405
box -295 -319 295 319
use sky130_fd_pr__pfet_01v8_lvt_4Q3NH3  XM4
timestamp 1749567790
transform 1 0 2349 0 1 -1365
box -295 -319 295 319
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM6
timestamp 1749574077
transform 1 0 1321 0 1 -2186
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM7
timestamp 1749574077
transform 1 0 2343 0 1 -2186
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM8
timestamp 1749574077
transform 1 0 1329 0 1 -2962
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM9
timestamp 1749574077
transform 1 0 2359 0 1 -2966
box -211 -310 211 310
<< labels >>
flabel space 1558 68 1962 272 0 FreeSans 1600 0 0 0 Vdd
flabel space 564 -886 840 -746 0 FreeSans 480 0 0 0 Inn
flabel space 2798 -918 2932 -818 0 FreeSans 480 0 0 0 Inp
flabel space 2832 -3336 3080 -3236 0 FreeSans 480 0 0 0 Vss
flabel space 1014 -2620 1156 -2536 0 FreeSans 480 0 0 0 Ipn
flabel space 2490 -2594 2662 -2512 0 FreeSans 480 0 0 0 Ipp
flabel space 1634 -3630 1788 -3552 0 FreeSans 480 0 0 0 Vb2
flabel space 1998 -3628 2150 -3526 0 FreeSans 480 0 0 0 Vb3
flabel space 1342 -3648 1564 -3546 0 FreeSans 480 0 0 0 Vb1
flabel space 2780 -1862 3012 -1694 0 FreeSans 480 0 0 0 out
<< end >>
