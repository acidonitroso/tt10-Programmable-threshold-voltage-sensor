magic
tech sky130A
magscale 1 2
timestamp 1750067613
<< viali >>
rect -250 3800 -150 4100
rect -250 1300 -150 1600
rect -250 -1200 -150 -900
rect -250 -3750 -150 -3450
rect -250 -6350 -150 -6050
rect -250 -8700 -150 -8400
rect -250 -11350 -150 -11050
rect -250 -13700 -150 -13400
<< metal1 >>
rect -900 4100 -100 4150
rect -900 3800 -250 4100
rect -150 3800 -100 4100
rect -900 3750 -100 3800
rect -900 1650 -500 3750
rect -200 2050 100 3350
rect -900 1600 -100 1650
rect -900 1300 -250 1600
rect -150 1300 -100 1600
rect -900 1250 -100 1300
rect -900 -850 -500 1250
rect -200 -450 100 850
rect -900 -900 -100 -850
rect -900 -1200 -250 -900
rect -150 -1200 -100 -900
rect -900 -1250 -100 -1200
rect -900 -3400 -500 -1250
rect -200 -2950 100 -1650
rect -900 -3450 -100 -3400
rect -900 -3750 -250 -3450
rect -150 -3750 -100 -3450
rect -900 -3800 -100 -3750
rect -900 -6000 -500 -3800
rect -200 -5450 100 -4150
rect -900 -6050 -50 -6000
rect -900 -6350 -250 -6050
rect -150 -6350 -50 -6050
rect -900 -6400 -50 -6350
rect -900 -8350 -500 -6400
rect -200 -7950 100 -6650
rect -900 -8400 -100 -8350
rect -900 -8700 -250 -8400
rect -150 -8700 -100 -8400
rect -900 -8750 -100 -8700
rect -900 -11000 -500 -8750
rect -200 -10450 100 -9150
rect -900 -11050 -100 -11000
rect -900 -11350 -250 -11050
rect -150 -11350 -100 -11050
rect -900 -11400 -100 -11350
rect -900 -13350 -500 -11400
rect -200 -12950 100 -11650
rect -900 -13400 -100 -13350
rect -900 -13700 -250 -13400
rect -150 -13700 -100 -13400
rect -900 -13750 -100 -13700
use sky130_fd_pr__res_high_po_0p35_3S7HW9  sky130_fd_pr__res_high_po_0p35_3S7HW9_0
timestamp 1750063742
transform 1 0 -49 0 1 -11038
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  sky130_fd_pr__res_high_po_0p35_3S7HW9_2
timestamp 1750063742
transform 1 0 -49 0 1 3962
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  sky130_fd_pr__res_high_po_0p35_3S7HW9_3
timestamp 1750063742
transform 1 0 -49 0 1 1462
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  XR14
timestamp 1750063742
transform 1 0 -49 0 1 -1038
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  XR15
timestamp 1750063742
transform 1 0 -49 0 1 -3538
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  XR16
timestamp 1750063742
transform 1 0 -49 0 1 -6038
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  XR17
timestamp 1750063742
transform 1 0 -49 0 1 -8538
box -201 -1212 201 1212
use sky130_fd_pr__res_high_po_0p35_3S7HW9  XR18
timestamp 1750063742
transform 1 0 -49 0 1 -13538
box -201 -1212 201 1212
<< end >>
