magic
tech sky130A
magscale 1 2
timestamp 1749574077
<< error_p >>
rect -223 181 -161 187
rect -95 181 -33 187
rect 33 181 95 187
rect 161 181 223 187
rect -223 147 -211 181
rect -95 147 -83 181
rect 33 147 45 181
rect 161 147 173 181
rect -223 141 -161 147
rect -95 141 -33 147
rect 33 141 95 147
rect 161 141 223 147
rect -223 -147 -161 -141
rect -95 -147 -33 -141
rect 33 -147 95 -141
rect 161 -147 223 -141
rect -223 -181 -211 -147
rect -95 -181 -83 -147
rect 33 -181 45 -147
rect 161 -181 173 -147
rect -223 -187 -161 -181
rect -95 -187 -33 -181
rect 33 -187 95 -181
rect 161 -187 223 -181
<< nwell >>
rect -423 -319 423 319
<< pmoslvt >>
rect -227 -100 -157 100
rect -99 -100 -29 100
rect 29 -100 99 100
rect 157 -100 227 100
<< pdiff >>
rect -285 88 -227 100
rect -285 -88 -273 88
rect -239 -88 -227 88
rect -285 -100 -227 -88
rect -157 88 -99 100
rect -157 -88 -145 88
rect -111 -88 -99 88
rect -157 -100 -99 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 99 88 157 100
rect 99 -88 111 88
rect 145 -88 157 88
rect 99 -100 157 -88
rect 227 88 285 100
rect 227 -88 239 88
rect 273 -88 285 88
rect 227 -100 285 -88
<< pdiffc >>
rect -273 -88 -239 88
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect 239 -88 273 88
<< nsubdiff >>
rect -387 249 -291 283
rect 291 249 387 283
rect -387 187 -353 249
rect 353 187 387 249
rect -387 -249 -353 -187
rect 353 -249 387 -187
rect -387 -283 -291 -249
rect 291 -283 387 -249
<< nsubdiffcont >>
rect -291 249 291 283
rect -387 -187 -353 187
rect 353 -187 387 187
rect -291 -283 291 -249
<< poly >>
rect -227 181 -157 197
rect -227 147 -211 181
rect -173 147 -157 181
rect -227 100 -157 147
rect -99 181 -29 197
rect -99 147 -83 181
rect -45 147 -29 181
rect -99 100 -29 147
rect 29 181 99 197
rect 29 147 45 181
rect 83 147 99 181
rect 29 100 99 147
rect 157 181 227 197
rect 157 147 173 181
rect 211 147 227 181
rect 157 100 227 147
rect -227 -147 -157 -100
rect -227 -181 -211 -147
rect -173 -181 -157 -147
rect -227 -197 -157 -181
rect -99 -147 -29 -100
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect -99 -197 -29 -181
rect 29 -147 99 -100
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 29 -197 99 -181
rect 157 -147 227 -100
rect 157 -181 173 -147
rect 211 -181 227 -147
rect 157 -197 227 -181
<< polycont >>
rect -211 147 -173 181
rect -83 147 -45 181
rect 45 147 83 181
rect 173 147 211 181
rect -211 -181 -173 -147
rect -83 -181 -45 -147
rect 45 -181 83 -147
rect 173 -181 211 -147
<< locali >>
rect -387 249 -291 283
rect 291 249 387 283
rect -387 187 -353 249
rect 353 187 387 249
rect -227 147 -211 181
rect -173 147 -157 181
rect -99 147 -83 181
rect -45 147 -29 181
rect 29 147 45 181
rect 83 147 99 181
rect 157 147 173 181
rect 211 147 227 181
rect -273 88 -239 104
rect -273 -104 -239 -88
rect -145 88 -111 104
rect -145 -104 -111 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 111 88 145 104
rect 111 -104 145 -88
rect 239 88 273 104
rect 239 -104 273 -88
rect -227 -181 -211 -147
rect -173 -181 -157 -147
rect -99 -181 -83 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 83 -181 99 -147
rect 157 -181 173 -147
rect 211 -181 227 -147
rect -387 -249 -353 -187
rect 353 -249 387 -187
rect -387 -283 -291 -249
rect 291 -283 387 -249
<< viali >>
rect -211 147 -173 181
rect -83 147 -45 181
rect 45 147 83 181
rect 173 147 211 181
rect -273 -88 -239 88
rect -145 -88 -111 88
rect -17 -88 17 88
rect 111 -88 145 88
rect 239 -88 273 88
rect -211 -181 -173 -147
rect -83 -181 -45 -147
rect 45 -181 83 -147
rect 173 -181 211 -147
<< metal1 >>
rect -223 181 -161 187
rect -223 147 -211 181
rect -173 147 -161 181
rect -223 141 -161 147
rect -95 181 -33 187
rect -95 147 -83 181
rect -45 147 -33 181
rect -95 141 -33 147
rect 33 181 95 187
rect 33 147 45 181
rect 83 147 95 181
rect 33 141 95 147
rect 161 181 223 187
rect 161 147 173 181
rect 211 147 223 181
rect 161 141 223 147
rect -279 88 -233 100
rect -279 -88 -273 88
rect -239 -88 -233 88
rect -279 -100 -233 -88
rect -151 88 -105 100
rect -151 -88 -145 88
rect -111 -88 -105 88
rect -151 -100 -105 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 105 88 151 100
rect 105 -88 111 88
rect 145 -88 151 88
rect 105 -100 151 -88
rect 233 88 279 100
rect 233 -88 239 88
rect 273 -88 279 88
rect 233 -100 279 -88
rect -223 -147 -161 -141
rect -223 -181 -211 -147
rect -173 -181 -161 -147
rect -223 -187 -161 -181
rect -95 -147 -33 -141
rect -95 -181 -83 -147
rect -45 -181 -33 -147
rect -95 -187 -33 -181
rect 33 -147 95 -141
rect 33 -181 45 -147
rect 83 -181 95 -147
rect 33 -187 95 -181
rect 161 -147 223 -141
rect 161 -181 173 -147
rect 211 -181 223 -147
rect 161 -187 223 -181
<< properties >>
string FIXED_BBOX -370 -266 370 266
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 0.35 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
