magic
tech sky130A
magscale 1 2
timestamp 1750071538
<< viali >>
rect 266 3600 336 3798
rect 832 3616 902 3814
<< metal1 >>
rect 76 6136 1098 6596
rect 246 3814 932 3822
rect 246 3798 832 3814
rect 246 3600 266 3798
rect 336 3616 832 3798
rect 902 3616 932 3814
rect 336 3600 932 3616
rect 246 3592 932 3600
rect 492 1917 706 3592
rect 854 1917 1188 2118
rect 492 1703 1188 1917
rect -394 1598 -196 1604
rect -394 1154 -196 1400
rect 854 1455 1188 1703
rect -398 694 208 1154
rect 854 1115 1188 1121
<< via1 >>
rect -394 1400 -196 1598
rect 854 1121 1188 1455
<< metal2 >>
rect -394 1819 -196 1828
rect -394 1598 -196 1621
rect -400 1400 -394 1598
rect -196 1400 -190 1598
rect 848 1121 854 1455
rect 1188 1121 1194 1455
rect 854 902 1188 911
<< via2 >>
rect -394 1621 -196 1819
rect 854 1121 1188 1245
rect 854 911 1188 1121
<< metal3 >>
rect -394 2025 -196 2031
rect -394 1824 -196 1827
rect -399 1819 -191 1824
rect -399 1621 -394 1819
rect -196 1621 -191 1819
rect -399 1616 -191 1621
rect 849 1245 1193 1250
rect 849 906 854 1245
rect 1188 906 1193 1245
rect 854 691 1188 697
<< via3 >>
rect -394 1827 -196 2025
rect 854 911 1188 1031
rect 854 697 1188 911
<< metal4 >>
rect -394 2026 -195 6601
rect -395 2025 -195 2026
rect -395 1827 -394 2025
rect -196 1827 -195 2025
rect -395 1826 -195 1827
rect 853 1031 1189 1032
rect 853 697 854 1031
rect 1188 697 1189 1031
rect 853 696 1189 697
rect 854 499 1188 696
use sky130_fd_pr__res_high_po_0p35_MGTKQ5  XR7 ~/tt10-analog-template-psei-def/mag
timestamp 1749664143
transform 1 0 148 0 1 3649
box -201 -3102 201 3102
use sky130_fd_pr__res_high_po_0p35_KC2364  XR8
timestamp 1749664143
transform 1 0 1017 0 1 4134
box -201 -2612 201 2612
<< labels >>
flabel space 316 6774 738 6970 0 FreeSans 1600 0 0 0 Vmirpmos
flabel space 1050 1208 1614 1598 0 FreeSans 1600 0 0 0 Vss
flabel space -918 6882 -228 7220 0 FreeSans 1600 0 0 0 Vdd
<< end >>
